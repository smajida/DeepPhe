|patient ID|cancer  link|body location|document for body location |body location clockface position|documents for body location clockface position|body location quadrant|documents for body location quadrant|clinical T classification|clinical N classification|clinical M classification|clinical prefix|clinical suffix|pathologic T classification|pathologic N classification|pathologic M classification|pathologic prefix|pathologic suffix|generic T classification|generic N classification|generic M classification|generic prefix|generic suffix|Diagnosis|document for diagnosis|tumor type|documents for tumor type|cancer type|documents for cancer type|histologic type|documents for histologic type|tumor extent|documents for extent|er status interpretation|documents for er status interpretation|er status numeric value|documents for er numeric value|er status method|documents for er status method|pr status interpretation|documents for pr status interpretation|pr status numeric value|documents for pr numeric value|pr status method|documents for pr status method|her2neu status interpretation|documents for her2neu status interpretation|her2neu status numeric value|documents for her2neu status numeric value|her2neu status method|documents for her2 status method
|patient04|cancer_13_patient04|Left_Breast|report002_RAD; report005_SP; report006_RAD; report008_RAD|1 o'clock position|report002_RAD; report005_SP; report006_RAD; report008_RAD;|Upper-Outer Quadrant of the Breast|report002_RAD; report006_RAD; report008_RAD||||||||||||||||Invasive_Lobular_Breast_Carcinoma; 
Lobular_Breast_Carcinoma_In_Situ|report005_SP; report006_RAD; report008_RAD|primary||Carcinoma||Lobular||In-Situ; 
Invasive||Positive|report005_SP|200|report005_SP|IHC|report005_SP|Positive|report005_SP|270|report005_SP|IHC|report005_SP|Negative|report005_SP|1+|report005_SP|IHC|report005_SP
