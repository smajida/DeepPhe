cancer ID|patient ID|body location|documents for|clinical stage|documents for clinical stage|clinical T classification|documents for clinical T classification|clinical N classification|documents for clinical N classification|clinical M classification|documents for clinical M classification|clinical prefix|documents for clinical prefix|clinical suffix|documents for clinical suffix|pathologic T classification|documents for pathologic T classification|pathologic N classification|documents for pathologic N classification|pathologic M classification|documents for pathologic M classification|pathologic prefix|documents for pathologic prefix|pathologic suffix|documents for pathologic suffix|generic T classification|documents for generic T classification|generic N classification|documents for generic N classification|generic M classification|documents for generic M classification|generic prefix|documents for generic prefix|generic suffix|documents for generic suffix
cancer_12_patient04|patient04|Left_Breast|report002_RAD; report005_SP; report008_RAD||||||||||||||||||||||||||||||||
