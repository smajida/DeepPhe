C0524811|T061|Fractionation
C0524811|T061|Radiotherapy Dose Fractionations
C0524811|T061|Dose Fractionations
C0524811|T061|Fractionation, Dose
C0524811|T061|fractionation
C0524811|T061|Fractionation Radiotherapy
C0524811|T061|Dose Fractionation, Radiotherapy
C0524811|T061|Fractionations, Radiotherapy Dose
C0524811|T061|Fractionations, Dose
C0524811|T061|RADIOTHER DOSE FRACTIONATION
C0524811|T061|Fractionation, Radiotherapy Dose
C0524811|T061|Radiotherapy Dose Fractionation
C0524811|T061|Dose Fractionation
C0524811|T061|Dose Fractionations, Radiotherapy
C1335378|T191|Pericardial Carcinomatosis
C1335378|T191|Carcinomatosis of the Pericardium
C0456908|T033|N1b Stage Finding
C0456908|T033|N1b TNM Finding
C0456908|T033|N1b Stage
C0456908|T033|Lymph Node Stage N1b
C0456908|T033|N1b Lymph Node Stage
C0456908|T033|N1b Cancer Stage Finding
C0456908|T033|Node Stage N1b
C0456908|T033|N1b
C0456908|T033|Node stage N1b
C0456908|T033|N1b Lymph Node Finding
C0456908|T033|N1b Regional Lymph Nodes Finding
C0456908|T033|N1b Node Finding
C0456908|T033|Node stage N1b (finding)
C0456908|T033|N1b Regional Lymph Node Stage Finding
C0456908|T033|N1b Node Stage
C1514710|T061|High-LET Radiotherapy
C1514710|T061|high-dose radiation
C1514710|T061|Radiotherapy-High LET
C1514710|T061|Radiotherapy, High Linear Energy Transfer
C0855104|T191|Recurrent Burkitt Lymphoma
C0855104|T191|Relapsed Burkitt's Lymphoma
C0855104|T191|Recurrent Burkitt's Lymphoma
C0855104|T191|Burkitt's lymphoma recurrent
C0855104|T191|Burkitt's tumor or lymphoma recurrent
C0855104|T191|Burkitt's tumor recurrent
C0855104|T191|Burkitt's tumour recurrent
C0855104|T191|Burkitt's tumour or lymphoma recurrent
C0854839|T191|Recurrent Angioimmunoblastic T-cell Lymphoma
C0854839|T191|Relapsed Angioimmunoblastic T-cell Lymphoma
C0935909|T191|Breast Carcinoma Metastatic to the Skin
C0935909|T191|Cutaneous Breast Cancer
C0935909|T191|cutaneous breast cancer
C0278689|T191|Recurrent Ovarian Carcinoma
C0278689|T191|Ovarian cancer recurrent
C0278689|T191|ovarian cancer, recurrent
C0278689|T191|recurrent ovarian carcinoma
C0278689|T191|Recurrent Ovarian Epithelial Cancer
C0278689|T191|Recurrent Carcinoma of the Ovary
C0278689|T191|Relapsed Ovarian Carcinoma
C0278689|T191|Ovarian epithelial cancer recurrent
C0278689|T191|ovary cancer, recurrent
C0278689|T191|Recurrent Ovarian Cancer
C0278689|T191|Relapsed Carcinoma of Ovary
C0278689|T191|Recurrent Carcinoma of Ovary
C0278689|T191|Recurrent Epithelial Cancer of Ovary
C0278689|T191|Relapsed Ovarian Epithelial Cancer
C0278689|T191|recurrent ovarian epithelial cancer
C0278689|T191|Recurrent Epithelial Cancer of the Ovary
C0278689|T191|ovarian carcinoma, recurrent
C0278689|T191|recurrent ovary cancer
C0278689|T191|Relapsed Epithelial Cancer of Ovary
C0278689|T191|Relapsed Carcinoma of the Ovary
C0278689|T191|Relapsed Epithelial Cancer of the Ovary
C0278689|T191|ovarian epithelial cancer, recurrent
C0278689|T191|recurrent ovarian cancer
C1332986|T191|Childhood Osteosarcoma
C1332986|T191|Pediatric Osteosarcoma
C0007112|T191|Prostate Adenocarcinoma
C0007112|T191|PROSTATE, ADENOCARCINOMA
C0007112|T191|adenocarcinoma of the prostate
C0007112|T191|Adenocarcinoma of prostate (disorder)
C0007112|T191|prostate cancer, adenocarcinoma
C0007112|T191|Adenocarcinoma of Prostate
C0007112|T191|Adenocarcinoma of prostate
C0007112|T191|Adenocarcinoma of the Prostate
C0007112|T191|adenocarcinoma, prostatic
C0007112|T191|prostatic adenocarcinoma
C1883632|T045|3' Flank Mutation
C0577018|T033|Stomach Mass
C0577018|T033|Stomach mass
C0577018|T033|Mass of Stomach
C0577018|T033|Mass of the Stomach
C0577018|T033|Mass of stomach (finding)
C0577018|T033|Gastric Mass
C0577018|T033|Lump stomach
C0577018|T033|Mass of stomach
C0278580|T191|Recurrent Cutaneous T-Cell Non-Hodgkin Lymphoma
C0278580|T191|Recurrent Skin T-Cell Lymphoma
C0278580|T191|Recurrent Cutaneous T-Cell Non-Hodgkin's Lymphoma
C0278580|T191|Relapsed T-Cell Lymphoma of the Skin
C0278580|T191|Recurrent T-Cell Lymphoma of Skin
C0278580|T191|Relapsed T-Cell Lymphoma of Skin
C0278580|T191|Relapsed Skin T-Cell Lymphoma
C0278580|T191|Relapsed Cutaneous T-Cell Lymphoma
C0278580|T191|Recurrent T-Cell Lymphoma of the Skin
C0278787|T191|Recurrent Chronic Myelogenous Leukemia, BCR-ABL1 Positive
C0278787|T191|Recurrent Chronic Myelogenous Leukemia
C0278787|T191|Relapsed CML
C0278787|T191|Relapsed Chronic Myelogenous Leukemia
C0278787|T191|Relapsed CGL
C1883643|T045|5' Flank Mutation
C0855042|T191|Metastatic Extraosseous Ewing Sarcoma
C0855042|T191|Extra-Osseous Ewing's Sarcoma, Metastatic
C0855042|T191|Metastatic Extra-Osseous Ewing's Sarcoma
C0855042|T191|Extra-osseous Ewing's sarcoma metastatic
C0855042|T191|Metastatic Extraskeletal Ewing's Sarcoma
C0855042|T191|Metastatic Extraosseous Ewing's Sarcoma
C2347442|T033|Palisading Necrosis
C0855050|T191|Metastatic Extraskeletal Osteosarcoma
C0855050|T191|Extraskeletal Osteosarcoma, Metastatic
C0855050|T191|Extraskeletal osteosarcoma metastatic
C0855050|T191|Metastatic Extraosseous Osteosarcoma
C0855050|T191|Metastatic Extraskeletal Osteogenic Sarcoma
C1332050|T191|AIDS-Related Malignant Cervical Neoplasm
C1332050|T191|AIDS-Related Malignant Neoplasm of the Cervix Uteri
C1332050|T191|AIDS-Related Malignant Neoplasm of Uterine Cervix
C1332050|T191|AIDS-Related Malignant Neoplasm of Cervix
C1332050|T191|AIDS-Related Malignant Cervix Uteri Neoplasm
C1332050|T191|AIDS-Related Malignant Cervix Neoplasm
C1332050|T191|AIDS-Related Malignant Neoplasm of the Cervix
C1332050|T191|AIDS-Related Malignant Neoplasm of Cervix Uteri
C1332050|T191|AIDS-Related Malignant Cervix Tumor
C1332050|T191|AIDS-Related Malignant Cervical Tumor
C1332050|T191|AIDS-Related Malignant Tumor of the Cervix Uteri
C1332050|T191|AIDS-Related Malignant Tumor of the Uterine Cervix
C1332050|T191|AIDS-Related Malignant Tumor of Cervix
C1332050|T191|AIDS-Related Malignant Uterine Cervix Neoplasm
C1332050|T191|AIDS-Related Malignant Uterine Cervix Tumor
C1332050|T191|AIDS-Related Malignant Tumor of Uterine Cervix
C1332050|T191|AIDS-Related Malignant Cervix Uteri Tumor
C1332050|T191|AIDS-Related Malignant Tumor of Cervix Uteri
C1332050|T191|AIDS-Related Malignant Tumor of the Cervix
C1332050|T191|AIDS-Related Malignant Neoplasm of the Uterine Cervix
C0024884|T061|Radical Mastectomy
C0024884|T061|Halsted radical mastectomy
C0024884|T061|Mastectomies, Radical
C0024884|T061|Radical mastectomy (procedure)
C0024884|T061|Mastectomy, Radical
C0024884|T061|Mastectomy radical
C0024884|T061|RADICAL MASTECTOMY
C0024884|T061|Radical Mastectomies
C0024884|T061|Radical mastectomy including pectoral muscles and axillary lymph nodes
C0024884|T061|radical mastectomy
C0024884|T061|Halsted Radical Mastectomy
C0024884|T061|Radical mastectomy including pectoral muscles and axillary lymph nodes (procedure)
C0024884|T061|Radical mastectomy NOS
C0024884|T061|Radical mastectomy
C0686114|T191|Metastatic Malignant Neoplasm to the Extrahepatic Bile Ducts
C1333012|T191|Childhood Testicular Yolk Sac Tumor
C1333012|T191|Childhood Testicular Yolk Sac Neoplasm
C1333012|T191|Pediatric Testicular Endodermal Sinus Tumor
C1333012|T191|Childhood Testicular Endodermal Sinus Tumor
C1333012|T191|Childhood Testicular Endodermal Sinus Neoplasm
C1333012|T191|Pediatric Testicular Yolk Sac Neoplasm
C1333012|T191|Pediatric Testicular Endodermal Sinus Neoplasm
C1333012|T191|Pediatric Testicular Yolk Sac Tumor
C2987252|T191|Esophageal Spindle Cell Carcinoma
C2987252|T191|Esophageal Carcinoma with Mesenchymal Stroma
C2987252|T191|Esophageal Pseudosarcomatous Squamous Cell Carcinoma
C2987252|T191|Esophageal Carcinosarcoma
C2987252|T191|Esophageal Squamous Cell Carcinoma with a Spindle-Cell Component
C2987252|T191|Esophageal Sarcomatoid Carcinoma
C2987252|T191|Esophageal Metaplastic Carcinoma
C2987252|T191|Esophageal Polypoid Carcinoma
C1513784|T061|Myeloablative Chemotherapy
C1513784|T061|myeloablative chemotherapy
C3179062|T061|Image Guided Radiation Therapy
C3179062|T061|IGRT
C3179062|T061|Radiation Therapies, Image-Guided
C3179062|T061|Radiation Therapy, Image-Guided
C3179062|T061|Radiotherapy, Image Guided
C3179062|T061|Radiotherapies, Image-Guided
C3179062|T061|Therapies, Image-Guided Radiation
C3179062|T061|Radiotherapy, Image-Guided
C3179062|T061|image-guided radiation therapy
C3179062|T061|Therapy, Image-Guided Radiation
C3179062|T061|Image-Guided Radiation Therapies
C3179062|T061|Image-Guided Radiotherapy
C3179062|T061|Image-Guided Radiation Therapy
C3179062|T061|Image-Guided Radiotherapies
C1335705|T191|Recurrent Male Reproductive System Carcinoma
C1335705|T191|Recurrent Male Reproductive System Cancer
C0544886|T049|Somatic Mutation
C0544886|T049|Somatic Mutation Abnormality
C0544886|T049|Somatic mutation (finding)
C0544886|T049|somatic mutation
C0544886|T049|Somatic mutation
C0475394|T185|T3c Stage Finding
C0475394|T185|Tumor Stage T3c
C0475394|T185|T3c tumor stage
C0475394|T185|T3c Primary Tumor Stage Finding
C0475394|T185|Tumour stage T3c
C0475394|T185|T3c Primary Tumor Finding
C0475394|T185|T3c Stage
C0475394|T185|Tumor stage T3c (finding)
C0475394|T185|T3c Cancer Stage Finding
C0475394|T185|T3c Tumor Finding
C0475394|T185|T3c
C0475394|T185|T3c TNM Finding
C0475394|T185|Tumor stage T3c
C0475394|T185|T3c Tumor Stage
C0475387|T185|T2a Stage Finding
C0475387|T185|T2a Cancer Stage Finding
C0475387|T185|T2a Tumor Stage
C0475387|T185|T2a TNM Finding
C0475387|T185|T2a Stage
C0475387|T185|Tumour stage T2a
C0475387|T185|T2a Tumor Finding
C0475387|T185|Tumor Stage T2a
C0475387|T185|T2a Primary Tumor Stage Finding
C0475387|T185|T2a
C0475387|T185|Tumor stage T2a (finding)
C0475387|T185|T2a Primary Tumor Finding
C0475387|T185|Tumor stage T2a
C1522058|T046|Coagulative Necrosis
C1522058|T046|Coagulative necrosis
C1522058|T046|Coagulative necrosis (morphologic abnormality)
C1522058|T046|Coagulation necrosis
C1336735|T191|Therapy-Related Acute Myeloid Leukemia
C1336735|T191|Treatment-Related AML
C1336735|T191|Treatment related acute myeloid leukemia
C1336735|T191|Treatment related AML
C1336735|T191|Treatment-related Acute Myeloid Leukemia
C1336735|T191|Treatment-Related Acute Myelocytic Leukemia
C1336735|T191|Treatment Related Acute Myelocytic Leukemia
C1336735|T191|Treatment Related Acute Myeloid Leukemia
C1336735|T191|Treatment Related Acute Myelogenous Leukemia
C1336735|T191|t-AML
C1336735|T191|Treatment Related AML
C1336735|T191|Treatment-Related Acute Myelogenous Leukemia
C0278775|T191|Recurrent Adult Liver Carcinoma
C0278775|T191|Relapsed Adult Liver Cancer
C0278775|T191|Relapsed Adult Primary Liver Cancer
C0278775|T191|hepatoma, recurrent adult primary
C0278775|T191|Relapsed Adult Primary Cancer of Liver
C0278775|T191|Recurrent Adult Primary Cancer of Liver
C0278775|T191|recurrent adult primary liver cancer
C0278775|T191|adult primary hepatoma, recurrent
C0278775|T191|Recurrent Adult Primary Liver Cancer
C0278775|T191|Recurrent Adult Liver Cancer
C0278775|T191|liver cancer, recurrent adult primary
C0278775|T191|adult primary liver cancer, recurrent
C0278775|T191|Recurrent Adult Primary Cancer of the Liver
C0278775|T191|Relapsed Adult Primary Cancer of the Liver
C1332284|T191|Anaplastic Lymphoma Post-Transplant Lymphoproliferative Disorder
C1332284|T191|Anaplastic Diffuse Large B-Cell Lymphoma PTLD
C1332284|T191|Anaplastic Lymphoma PTLD
C0854825|T191|Stage IV Anaplastic Large Cell Lymphoma
C0854825|T191|Anaplastic Large Cell Lymphoma T- and Null-Cell Types Stage IV
C0854825|T191|Anaplastic Large Cell Lymphoma Stage IV
C0246421|T121|Letrozole
C0246421|T121|letrozole
C0246421|T121|LETROZOLE
C0246421|T121|4,4'-(1H-1,2,4triazol-1-ylmethylene)dibenzonitrile
C0246421|T121|CGS 20267
C0246421|T121|Femara
C0195495|T061|Bilateral Salpingectomy with Oophorectomy
C0195495|T061|bilateral salpingo-oophorectomy
C0341353|T047|Appendix Mass
C0341353|T047|Appendix mass
C0341353|T047|Mass of appendix (finding)
C0341353|T047|Appendiceal Mass
C0341353|T047|Mass of appendix
CL388688|T191|Sarcomatoid Squamous Cell Carcinoma
CL388688|T191|Spindle Cell (Sarcomatoid) Squamous Cell Carcinoma
CL388688|T191|Epidermoid carcinoma - spindle cell
CL388688|T191|Squamous cell carcinoma - spindle cell
CL388688|T191|Epidermoid carcinoma, spindle cell
CL388688|T191|Squamous cell carcinoma, spindle cell
CL388688|T191|Squamous cell carcinoma, sarcomatoid
CL388688|T191|Squamous Cell Carcinoma, Spindle Cell
CL388688|T191|Squamous Cell Spindle Cell Carcinoma
CL388688|T191|Spindle cell squamous cell carcinoma (disorder)
CL388688|T191|Epidermoid Spindle Cell Carcinoma
CL388688|T191|Spindle cell squamous cell carcinoma
CL388688|T191|Squamous cell carcinoma, spindle cell (morphologic abnormality)
CL388688|T191|Squamous Cell Carcinoma, Sarcomatoid
C1301095|T201|Size of base of tumor on transillumination
C1301095|T201|Size of base of tumor on transillumination (observable entity)
C1301095|T201|Size of base of tumour on transillumination
C0333514|T046|Zonal Necrosis
C0333514|T046|Zonal necrosis
C0333514|T046|Zonal necrosis (morphologic abnormality)
C2986463|T034|Androgen Receptor Positive
C2986463|T034|AR+
C2986463|T034|androgen receptor positive
C1335663|T033|Rapidly Enlarging Mass
C0449453|T082|Lesion size
C0449453|T082|Size of lesion
C0449453|T082|Lesion size (observable entity)
C1334786|T191|Mixed Hepatoblastoma with Teratoid Features
C1332624|T191|Breast Carcinoma Metastatic to the Brain
C0449455|T082|Calculus size
C0449455|T082|Size of calculus
C0449455|T082|Calculus size (observable entity)
C1336869|T191|Unresectable Malignant Neoplasm
C1336869|T191|Unresectable Malignant Tumor
C0854824|T191|Stage III Anaplastic Large Cell Lymphoma
C0854824|T191|Anaplastic Large Cell Lymphoma Stage III
C0854824|T191|Anaplastic Large Cell Lymphoma T- and Null-Cell Types Stage III
C0349543|T191|Brain Glioblastoma
C0349543|T191|Grade IV Brain Astrocytic Tumor
C0349543|T191|Grade IV Astrocytic Neoplasm of Brain
C0349543|T191|Grade IV Astrocytic Neoplasm of the Brain
C0349543|T191|Grade IV Brain Astrocytic Neoplasm
C0349543|T191|Glioblastoma multiforme of brain
C0349543|T191|Glioblastoma multiforme of brain (disorder)
C0349543|T191|Brain Glioblastoma Multiforme
C0349543|T191|Glioblastoma Multiforme of Brain
C0349543|T191|Grade IV Astrocytic Tumor of Brain
C0349543|T191|Glioblastoma Multiforme of the Brain
C0349543|T191|Grade IV Astrocytic Tumor of the Brain
C1334728|T191|Metastatic Malignant Neoplasm to the Iris
C1334728|T191|Metastatic Neoplasm to the Iris
C1334728|T191|Metastatic Tumor to the Iris
C0862402|T191|Stage II Bladder Urothelial Carcinoma
C0862402|T191|Stage II Urinary Bladder Transitional Cell Carcinoma
C0862402|T191|Stage II Bladder Urothelial Carcinoma AJCC v6
C0862402|T191|Stage II Bladder Urothelial Carcinoma AJCC v7
C0862402|T191|Stage II Transitional Cell Carcinoma of Bladder
C0862402|T191|Stage II Transitional Cell Carcinoma of the Bladder
C0862402|T191|Stage II Transitional Cell Carcinoma of Urinary Bladder
C0862402|T191|Stage II Transitional Cell Carcinoma of the Urinary Bladder
C3494227|T061|Craniospinal Irradiation
C3494227|T061|Spinocranial Irradiation
C3494227|T061|Irradiation, Spinocranial
C3494227|T061|craniospinal irradiation
C3494227|T061|Irradiation, Craniospinal
C3494227|T061|CSI
C1332626|T191|Breast Carcinoma Metastatic to the Lung
C1297883|T047|Radial Scar/Complex Sclerosing Lesion
C1297883|T047|Radial Scar
C1297883|T047|Radial Sclerosing Lesion
C1297883|T047|Complex Sclerosing Lesion
C1511316|T191|Breast Large Cell Neuroendocrine Carcinoma
C1300683|T074|CyberKnife
C1300683|T074|CyberKnife (physical object)
C0346957|T191|Disseminated Malignant Neoplasm
C0346957|T191|Generalized cancer
C0346957|T191|Disseminated cancer
C0346957|T191|Generalised cancer
C0346957|T191|CA - Disseminated cancer
C0346957|T191|Generalised malignancy
C0346957|T191|Disseminated malignancy
C0346957|T191|Widespread metastatic malignant neoplastic disease (disorder)
C0346957|T191|Malig neo disseminated
C0346957|T191|Disseminated malignant neoplasm without specification of site
C0346957|T191|Malignant neoplasm disseminated
C0346957|T191|Generalized malignancy
C0346957|T191|Disseminated malignant neoplasm
C0346957|T191|Widespread metastatic malignant neoplastic disease
C0346957|T191|Malignant neoplasm, disseminated
C1334279|T191|Invasive Micropapillary Breast Carcinoma
C1334279|T191|Infiltrating Micropapillary Breast Carcinoma
C0441905|T033|Venous stage VX
C0441905|T033|VX Venous Invasion Finding
C0441905|T033|VX: venous invasion cannot be assessed
C0441905|T033|VX stage (finding)
C0441905|T033|VX Stage Finding
C0441905|T033|VX TNM Finding
C0441905|T033|VX
C0441905|T033|Venous Stage VX
C0441905|T033|VX Stage
C0441905|T033|VX Cancer Stage Finding
C0441905|T033|VX Venous Stage
C0441905|T033|VX stage
C0346998|T191|Metastatic Malignant Neoplasm to the Vulva
C0346998|T191|Metastasis to the Vulva
C0346998|T191|Vulvar Metastasis
C0346998|T191|Metastatic Neoplasm to the Vulva
C1334928|T033|Necrotic Change
C1334928|T033|Necrotic changes (finding)
C1334928|T033|Necrotic changes
C1334928|T033|Necrosis
C1335255|T191|PRETEXT Stage 1 Hepatoblastoma
C0281702|T191|Stage II Childhood Burkitt Lymphoma
C0281702|T191|Stage II Childhood Small Non-Cleaved Cell Lymphoma
C0281702|T191|Stage II Pediatric Small Non-Cleaved Cell Lymphoma
C0281702|T191|Pediatric Small Non-Cleaved Cell Lymphoma Stage II
C0281702|T191|Childhood Small Non-Cleaved Cell Lymphoma Stage II
C0281702|T191|Stage II Childhood Burkitt's Lymphoma
C2348908|T034|HER2/Neu Negative
C2348908|T034|ERBB2 Negative
C1274073|T201|Tumor size, additional dimension
C1274073|T201|Tumour size, additional dimension
C1274073|T201|Tumor size, additional dimension (observable entity)
C0206180|T191|Systemic Anaplastic Large Cell Lymphoma
C0206180|T191|LYMPHOMA LARGE CELL KI 01
C0206180|T191|CD 030 POSITIVE ANAPLASTIC LARGE CELL LYMPHOMA
C0206180|T191|Lymphoma, Large-Cell, Anaplastic [Disease/Finding]
C0206180|T191|Anaplastic large cell lymphoma, systemic type
C0206180|T191|Systemic Anaplastic Large-Cell Lymphoma
C0206180|T191|Anaplastic large cell lymphoma T- and null-cell types
C0206180|T191|Anaplastic large cell lymphoma, CD30-positive
C0206180|T191|Anaplastic large-cell lymphoma, primary systemic type
C0206180|T191|Anaplastic large cell lymphoma, CD30+
C0206180|T191|Ki-1 Lymphoma
C0206180|T191|Anaplastic large cell lymphoma (ALCL) CD30+
C0206180|T191|anaplastic large cell lymphoma
C0206180|T191|Anaplastic large cell lymphoma, NOS
C0206180|T191|(Ki-1+) lymphoma
C0206180|T191|Large cell (Ki-1+) lymphoma [obs]
C0206180|T191|Anaplastic large cell lymphoma T- and null-cell types NOS
C0206180|T191|ANAPLASTIC LARGE CELL LYMPHOMA
C0206180|T191|Ki 1 Lymphoma
C0206180|T191|Large-Cell Lymphoma, Anaplastic
C0206180|T191|Ki-1+ ALCL
C0206180|T191|Anaplastic Large-Cell Lymphoma
C0206180|T191|CD30+ Anaplastic Large-Cell Lymphoma
C0206180|T191|Lymphoma, Anaplastic Large-Cell
C0206180|T191|Lymphoma, Large-Cell, Anaplastic
C0206180|T191|Large-Cell Lymphomas, Anaplastic
C0206180|T191|Ki-1 Lymphomas
C0206180|T191|Lymphomas, Ki-1
C0206180|T191|CD30 Positive Anaplastic Large Cell Lymphoma
C0206180|T191|Lymphoma, Large-Cell, Ki-1
C0206180|T191|lymphoma, anaplastic large cell
C0206180|T191|ALCL, systemic
C0206180|T191|Anaplastic large cell lymphoma
C0206180|T191|Anaplastic Large-Cell Lymphomas
C0206180|T191|Anaplastic large cell lymphomas T- and null-cell types
C0206180|T191|Anaplastic large-cell lymphoma
C0206180|T191|Large cell anaplastic lymphoma (disorder)
C0206180|T191|Ki-1+ Anaplastic Large Cell Lymphoma
C0206180|T191|ALCL
C0206180|T191|Large cell anaplastic lymphoma
C0206180|T191|CD30-Positive Anaplastic Large-Cell Lymphoma
C0206180|T191|Anaplastic Large Cell Lymphoma
C0206180|T191|CD30+ Anaplastic Large Cell Lymphoma
C0206180|T191|Lymphomas, Anaplastic Large-Cell
C0206180|T191|Lymphoma, Ki-1
C0206180|T191|Anaplastic large cell lymphoma, T cell and Null cell type (morphologic abnormality)
C0206180|T191|Anaplastic large cell lymphoma, T cell and Null cell type
C0854914|T191|Bilateral Retinoblastoma
C0854914|T191|Retinoblastoma bilateral
C1512747|T191|Infiltrating Bladder Urothelial Carcinoma with Glandular Differentiation
C1512747|T191|nfiltrating Bladder Urothelial Carcinoma with Glandular Differentiation
C1332994|T191|Childhood Parosteal Osteosarcoma
C1332994|T191|Childhood Parosteal Osteogenic Sarcoma
C0854959|T191|Recurrent Vulvar Carcinoma
C0854959|T191|carcinoma of the vulva, recurrent
C0854959|T191|Recurrent Vulvar Cancer
C0854959|T191|Relapsed Cancer of the Vulva
C0854959|T191|Vulval cancer recurrent
C0854959|T191|recurrent cancer of the vulva
C0854959|T191|Relapsed Vulvar Cancer
C0854959|T191|recurrent carcinoma of the vulva
C0854959|T191|Recurrent Cancer of Vulva
C0854959|T191|vulva cancer, recurrent
C0854959|T191|Relapsed Cancer of Vulva
C0854959|T191|cancer of the vulva, recurrent
C0854959|T191|vulvar cancer, recurrent
C0854959|T191|recurrent vulvar cancer
C0854959|T191|Recurrent Cancer of the Vulva
C0854959|T191|Relapsed Vulva Cancer
C0854959|T191|Recurrent Vulva Cancer
C0854959|T191|recurrent vulva cancer
C0685110|T191|Metastatic Malignant Neoplasm to the Heart
C0685110|T191|Metastatic Neoplasm to the Heart
C0685110|T191|Metastases to Heart
C0685110|T191|Metastasis to Heart
C0685110|T191|Metastatic Tumor to the Heart
C0685110|T191|Metastasis to the Heart
C0685110|T191|Metastases to the Heart
C1519487|T191|Squamous Cell Breast Carcinoma, Spindle Cell Variant
CL448373|T191|Recurrent Urethra Carcinoma
CL448373|T191|Relapsed Cancer of Urethra
CL448373|T191|Recurrent Cancer of the Urethra
CL448373|T191|Recurrent Urethra Cancer
CL448373|T191|urethral cancer, recurrent
CL448373|T191|Recurrent Cancer of Urethra
CL448373|T191|Relapsed Urethra Cancer
CL448373|T191|Relapsed Cancer of the Urethra
CL448373|T191|Recurrent Urethral Cancer
CL448373|T191|Relapsed Urethral Cancer
CL448373|T191|Relapsed Urethra Carcinoma
CL448373|T191|recurrent urethral cancer
CL448373|T191|Urethral Cancer, Recurrent
C0020632|T061|Hypophysectomy
C0020632|T061|Pituitectomy NOS
C0020632|T061|Excision of the Pituitary Gland
C0020632|T061|pituitectomy
C0020632|T061|Hypophysectomy NOS
C0020632|T061|Pituitectomy
C0020632|T061|Excision of the Pituitary Gland+B3297
C0020632|T061|Excision of pituitary gland
C0020632|T061|hypophysectomy
C0020632|T061|Hypophysectomies
C0020632|T061|Total excision of pituitary gland, unspecified approach
C0020632|T061|Hypophysis Excision
C0020632|T061|Excision of the Hypophysis
C0020632|T061|Hypophysis Cerebri Excision
C0020632|T061|Hypophysectomy (procedure)
C0020632|T061|Total exc pituitary NOS
C0020632|T061|Pituitary Gland Excision
C1706721|T061|Adjuvant Radiation Therapy
C0279985|T191|Childhood Alveolar Soft Part Sarcoma
C0279985|T191|sarcoma, alveolar soft-part, childhood
C0279985|T191|Pediatric Alveolar Soft Part Sarcoma
C0279985|T191|sarcoma, alveolar soft-part, pediatric
C0279985|T191|Childhood Alveolar Soft-Part Sarcoma
C0279985|T191|soft-part sarcoma, alveolar, childhood
C0279985|T191|soft-part sarcoma, alveolar, pediatric
C0279985|T191|childhood alveolar soft-part sarcoma
C0279985|T191|alveolar soft-part sarcoma, pediatric
C0279985|T191|alveolar soft-part sarcoma, childhood
C0279985|T191|pediatric alveolar soft-part sarcoma
C1335257|T191|PRETEXT Stage 3 Hepatoblastoma
C1883029|T191|Invasive Lobular Breast Carcinoma, Signet Ring Variant
C1883029|T191|Signet Ring Cell Lobular Breast Carcinoma
CL343405|T191|Recurrent Merkel Cell Carcinoma
CL343405|T191|recurrent neuroendocrine carcinoma of the skin
CL343405|T191|recurrent Merkel cell carcinoma
CL343405|T191|Merkel cell carcinoma, recurrent
CL343405|T191|Recurrent Neuroendocrine Carcinoma of the Skin
C0034619|T061|Radiation Therapy
C0034619|T061|Radiation
C0034619|T061|therapy, radiation
C0034619|T061|RADIOTHER
C0034619|T061|Therapeutic radiology
C0034619|T061|Therapeutic radiology procedure
C0034619|T061|irradiation
C0034619|T061|RADIATION
C0034619|T061|RADIATION THERAPY
C0034619|T061|Radiotherapy
C0034619|T061|Irradiation
C0034619|T061|RT
C0034619|T061|Radiation oncology AND/OR radiotherapy (procedure)
C0034619|T061|radiation therapy
C0034619|T061|Radiotherapy NOS
C0034619|T061|Irradiate
C0034619|T061|Radiotherapeutics
C0034619|T061|Radiation therapy
C0034619|T061|Radiation oncology AND/OR radiotherapy
C0034619|T061|Radiation Therapy Radiologic Technologist
C0034619|T061|radiotherapy
C0034619|T061|RT - Radiotherapy
C0034619|T061|Therapeutic radiology for cancer treatment
C0034619|T061|Irradiated
C0034619|T061|Therapy, Radiation
C0034619|T061|Cancer Radiotherapy
C0034619|T061|Radiotherapies
C0034619|T061|irradiated
C0334277|T191|Metastatic Adenocarcinoma
C0334277|T191|Adenocarcinoma, metastatic
C0334277|T191|Adenocarcinoma, metastatic (morphologic abnormality)
C0334277|T191|Adenocarcinoma, metastatic, NOS
C0334277|T191|Metastatic adenocarcinoma
C1370832|T191|Recurrent Childhood Hepatocellular Carcinoma
C1370832|T191|Recurrent Childhood Hepatoma
C1370832|T191|recurrent childhood hepatoma
C1370832|T191|hepatoma, pediatric, recurrent
C1370832|T191|Recurrent Pediatric Hepatoma
C1370832|T191|hepatoma, childhood, recurrent
C1370832|T191|pediatric hepatoma, recurrent
C1370832|T191|recurrent pediatric hepatoma
C1370832|T191|childhood hepatoma, recurrent
C1370832|T191|Recurrent Pediatric Hepatocellular Carcinoma
C0677984|T191|Locally Advanced Malignant Neoplasm
C0677984|T191|Locally Advanced Cancer
C0677984|T191|locally advanced cancer
C1883257|T061|TAC Regimen
C1883257|T061|Taxotere-Adriamycin-Cytoxan Regimen
C1883257|T061|TAC
C1883257|T061|Taxotere-Adriamycin-Cytoxan regimen
C1883257|T061|TAC regimen
C0184921|T060|Excisional Biopsy
C0184921|T060|surgical biopsy
C0184921|T060|Excisional biopsy
C0184921|T060|excisional biopsy
C0184921|T060|Excisional biopsy (procedure)
C0184921|T060|Excision biopsy (qualifier value)
C0184921|T060|Excision biopsy
CL447335|T061|Mini Ovoid Brachytherapy
C1333840|T191|Grade 2 Malignant Neoplasm
C115029|T191|Stage I Childhood Anaplastic Large Cell Lymphoma
C1515864|T191|Acinar Prostate Adenocarcinoma, Lymphoepithelioma-Like Variant
C120285|T081|Tumor Less Than or Equal to 2.0 Centimeters
C120285|T081|Less than or equal to 2.0 cm
C1516890|T049|Induced Gene Mutation
C1516890|T049|Environmentally Induced Gene Alteration
C1516890|T049|Environmentally Produced Alteration of Gene
C1516890|T049|Environmentally Produced Gene Alteration
C1516890|T049|Induced Gene Alteration
C1516890|T049|Gene Alteration, Environmentally Produced
C1516890|T049|Environmentally Induced Gene Mutation
C1709093|T049|Transition Mutation
C1709093|T049|Transition
C1709093|T049|Multiple Transition Abnormalities
C1709093|T049|transition mutation
C1709093|T049|Multiple Transition Mutations
C1709093|T049|Mutation, Transition
C1709093|T049|Transition Mutations
C1709093|T049|Nucleotide Transition Abnormality
C104990|T061|Retreatment of Progressive Local Disease with Brachytherapy
C0279915|T191|Stage I Childhood Hodgkin Lymphoma
C0279915|T191|Stage I Pediatric Hodgkin's Lymphoma
C0279915|T191|Childhood Hodgkin's Disease Stage I
C0279915|T191|Stage I Childhood Hodgkin's Lymphoma
C0279915|T191|Stage I Childhood Hodgkin's Disease
C0279915|T191|Pediatric Hodgkin's Lymphoma Stage I
C0279915|T191|Pediatric Hodgkin's Disease Stage I
C0279915|T191|stage I childhood Hodgkin lymphoma
C0279915|T191|Childhood Hodgkin's Lymphoma Stage I
C0279915|T191|Stage I Pediatric Hodgkin's Disease
C1333016|T191|Childhood Yolk Sac Tumor
C1333016|T191|Childhood Endodermal Sinus Neoplasm
C1333016|T191|Childhood Yolk Sac Neoplasm
C1333016|T191|Pediatric Endodermal Sinus Neoplasm
C1333016|T191|Childhood Endodermal Sinus Tumor
C1333016|T191|Pediatric Yolk Sac Tumor
C1333016|T191|Pediatric Yolk Sac Neoplasm
C1333985|T191|Hereditary Clear Cell Renal Cell Carcinoma
C1333985|T191|Hereditary Conventional (Clear Cell) Renal Cell Carcinoma
C2698204|T191|Metastatic Lobular Breast Carcinoma
C1336811|T191|Transplant-Related Hepatocellular Carcinoma
C1332942|T191|Childhood Anaplastic Large Cell Lymphoma
C1332942|T191|Pediatric CD30+ Anaplastic Large Cell Lymphoma
C1332942|T191|childhood anaplastic large cell lymphoma
C1332942|T191|Childhood K-1+ Anaplastic Large Cell Lymphoma
C1332942|T191|Childhood CD30+ Anaplastic Large Cell Lymphoma
C1332942|T191|Pediatric K-1+ Anaplastic Large Cell Lymphoma
C1332942|T191|Pediatric Anaplastic Large Cell Lymphoma
C111693|T191|Neural Glioblastoma
C0334459|T191|Infantile Fibrosarcoma
C0334459|T191|Congenital Fibrosarcoma
C0334459|T191|Infantile fibrosarcoma
C0334459|T191|Infantile fibrosarcoma (congenital fibrosarcoma)
C0334459|T191|Infantile fibrosarcoma (disorder)
C0334459|T191|Congenital fibrosarcoma
C0334459|T191|Infantile fibrosarcoma (morphologic abnormality)
C0024885|T061|Segmental Mastectomy
C0024885|T061|Segmental excision of breast (procedure)
C0024885|T061|Mastectomies, Segmental
C0024885|T061|Partial mastectomy (procedure)
C0024885|T061|Partial mastectomy
C0024885|T061|Mastectomies, Partial
C0024885|T061|Segmentectomy
C0024885|T061|Segmentectomies
C0024885|T061|Partial Mastectomy
C0024885|T061|segmental mastectomy
C0024885|T061|Partial Mastectomies
C0024885|T061|Mastectomy, Segmental
C0024885|T061|Subtotal mastectomy
C0024885|T061|Segmental excision of breast
C0024885|T061|Mastectomy, Partial
C0024885|T061|Excision of part of breast
C0024885|T061|PARTIAL MASTECTOMY
C0024885|T061|Segmental Mastectomies
C1708565|T191|Invasive Skin Melanoma
C1708565|T191|Infiltrating Melanoma
C1708565|T191|Invasive Melanoma
C0855111|T191|Recurrent Diffuse Large B-Cell Lymphoma
C0855111|T191|Relapsed Diffuse Large B-Cell Lymphoma
C2985436|T049|Deleterious Mutation
C2985436|T049|deleterious mutation
C3272465|T191|Ampulla of Vater Invasive Papillary Adenocarcinoma
C115363|T191|Recurrent Childhood Giant Cell Glioblastoma
C115363|T191|recurrent childhood giant cell glioblastoma
C0279069|T191|Recurrent Lymphomatoid Granulomatosis
C0279069|T191|Recurrent Angiocentric Immunoproliferative Lesion
C0279069|T191|Recurrent LYG
C0279069|T191|Relapsed Angiocentric Immunoproliferative Lesion
C1300096|T201|Tumor size, dimension 3
C1300096|T201|Tumour size, dimension 3
C1300096|T201|Tumor size, dimension 3 (observable entity)
C0475373|T033|T2 Stage Finding
C0475373|T033|T2 Stage
C0475373|T033|T2 Cancer Stage Finding
C0475373|T033|T2
C0475373|T033|Tumour stage T2
C0475373|T033|Tumor stage T2
C0475373|T033|T2 stage
C0475373|T033|T2 tumor stage
C0475373|T033|T2 Primary Tumor Finding
C0475373|T033|T2 category
C0475373|T033|T2 TNM Finding
C0475373|T033|T2 Tumor Stage
C0475373|T033|T2 Primary Tumor Stage Finding
C0475373|T033|T2 category (finding)
C0475373|T033|T2 Tumor Finding
C0475373|T033|Tumor Stage T2
C1300095|T201|Tumor size, dimension 2
C1300095|T201|Tumor size, dimension 2 (observable entity)
C1300095|T201|Tumour size, dimension 2
C1512920|T061|Intracavitary Radiation Therapy
C1512920|T061|Intracavitary Radiation
C1512920|T061|intracavitary radiation therapy
C0862643|T191|Stage IV Prostate Adenocarcinoma
C0862643|T191|Stage IV Prostate Adenocarcinoma AJCC v7
C1300094|T201|Tumor size, dimension 1
C1300094|T201|Tumor size, dimension 1 (observable entity)
C1300094|T201|Tumour size, dimension 1
C0279768|T034|Progesterone Receptor Status Unknown
C0279768|T034|unknown status, progesterone receptor
C0279768|T034|progesterone receptor status unknown
C0855153|T191|Recurrent Mediastinal (Thymic) Large B-Cell Cell Lymphoma
C0855153|T191|Relapsed Primary Mediastinal Large B-Cell Lymphoma
C0855153|T191|Recurrent Primary Mediastinal Large B-Cell Lymphoma
C0043162|T061|Total-Body Irradiation
C0043162|T061|Total Body Irradiation
C0043162|T061|TOTAL BODY IRRADIATION
C0043162|T061|Whole-Body Irradiation
C0043162|T061|total-body irradiation
C0195490|T061|Incomplete Oophorectomy
C0195490|T061|Partial excision of ovary
C0195490|T061|Partial oophorectomy
C0195490|T061|Incomplete Ovariectomy
C0195490|T061|Oophorectomy partial
C0195490|T061|Partial removal ovary
C0195490|T061|Ovariectomy, Incomplete
C0195490|T061|partial oophorectomy
C0195490|T061|Partial oophorectomy (procedure)
C0279561|T191|Tubular Breast Carcinoma
C0279561|T191|Infiltrating Tubular Carcinoma of Breast
C0279561|T191|tubular ductal breast carcinoma
C0279561|T191|Invasive Tubular Carcinoma of the Breast
C0279561|T191|Tubular breast carcinoma
C0279561|T191|Infiltrating Tubular Carcinoma of the Breast
C0279561|T191|Invasive Tubular Carcinoma of Breast
C0279561|T191|ductal tubular breast carcinoma
C0279561|T191|Invasive Tubular Breast Carcinoma
C0279561|T191|Infiltrating Tubular Breast Carcinoma
C0279561|T191|Tubular Carcinoma of Breast
C0279561|T191|Tubular Carcinoma of the Breast
C1720008|T191|AIDS-Related Burkitt Lymphoma
C1720008|T191|AIDS-Related Small Non-Cleaved Cell Lymphoma
C1720008|T191|AIDS Related Burkitt's Lymphoma
C1720008|T191|AIDS-Associated Burkitt's Lymphoma
C1720008|T191|AIDS-Associated Small Non Cleaved Cell Lymphoma
C1720008|T191|AIDS-Related Burkitt's Lymphoma
C1720008|T191|AIDS Related Small Non Cleaved Cell Lymphoma
CL472839|T191|Recurrent Combined Thymic Epithelial Neoplasm
C1516317|T033|Cauliflower-Like Mass
C0017636|T191|Glioblastoma
C0017636|T191|Glioblastoma, no ICD-O subtype
C0017636|T191|Glioblastoma, no ICD-O subtype (morphologic abnormality)
C0017636|T191|Glioblastomas
C0017636|T191|Grade IV Astrocytic Tumor
C0017636|T191|Astrocytomas, Grade IV
C0017636|T191|spongioblastoma multiforme
C0017636|T191|grade IV astrocytoma
C0017636|T191|Grade IV Astrocytic Neoplasm
C0017636|T191|GBM
C0017636|T191|BRAIN TUMOR, GLIOBLASTOMA MULTIFORME
C0017636|T191|Astrocytoma, Grade IV
C0017636|T191|Spongioblastoma Multiforme
C0017636|T191|Glioblastoma, NOS
C0017636|T191|Spongioblastoma multiforme
C0017636|T191|Glioblastoma multiforme
C0017636|T191|Glioblastoma Multiforme
C0017636|T191|Glioblastoma [Disease/Finding]
C0017636|T191|GLIOBLASTOMA MULTIFORME
C0017636|T191|astrocytoma WHO grade IV
C0017636|T191|GLM
C0017636|T191|glioblastoma
C0017636|T191|glioblastoma multiforme
C0017636|T191|SPONGIOBLASTOMA MULTIFORME
C0017636|T191|CANCER, GLIOBLASTOMA MULTIFORME
C0017636|T191|Grade IV Astrocytomas
C0017636|T191|INTRACRANIAL NEOPLASM, GLIOBLASTOMA MULTIFORME
C0017636|T191|Glioblastoma multiforme (disorder)
C0017636|T191|GBM - Glioblastoma multiforme
C0017636|T191|GLM - Glioblastoma multiforme
C0017636|T191|ASTROCYTOMA, GRADES 3-4
C0017636|T191|Grade IV Astrocytoma
C0017636|T191|GBM (Glioblastoma)
C1334704|T191|Metachronous Osteosarcoma
C1334704|T191|Metachronous Osteosarcoma of the Bone
C0424865|T033|Lump volume
C0424865|T033|Lump volume (observable entity)
C0424865|T033|Volume of lump
C0281704|T191|Stage III Childhood Burkitt Lymphoma
C0281704|T191|Stage III Pediatric Small Non-Cleaved Cell Lymphoma
C0281704|T191|Stage III Childhood Burkitt's Lymphoma
C0281704|T191|Childhood Small Non-Cleaved Cell Lymphoma Stage III
C0281704|T191|Stage III Childhood Small Non-Cleaved Cell Lymphoma
C0281704|T191|Pediatric Small Non-Cleaved Cell Lymphoma Stage III
C0279641|T191|Childhood Acute Promyelocytic Leukemia with t(15;17)(q22;q12); PML-RARA
C0279641|T191|M3 Childhood Acute Promyelocytic Leukemia
C0279641|T191|Childhood Acute Progranulocytic Leukemia
C0279641|T191|Childhood APL
C0279641|T191|Childhood Acute Promyelocytic Leukemia (M3)
C0279641|T191|Childhood M3 APL
C0279641|T191|Pediatric M3 APL
C0279641|T191|Pediatric Acute Promyelocytic Leukemia
C0279641|T191|Pediatric APL
C0279641|T191|M3 Pediatric Acute Promyelocytic Leukemia
C0279641|T191|Pediatric Acute M3 Leukemia
C0279641|T191|Pediatric Acute Progranulocytic Leukemia
C0279641|T191|Childhood Acute M3 Leukemia
C0279641|T191|Childhood Acute Promyelocytic Leukemia
C0454077|T061|Electron Beam Therapy
C0454077|T061|Teleradiotherapy using beta particles
C0454077|T061|electron beam therapy
C0454077|T061|Teleradiotherapy beta particles
C0454077|T061|photon beam radiation therapy
C0454077|T061|Electron teleradiotherap
C0454077|T061|Teleradiotherapy using electrons (procedure)
C0454077|T061|Betatron electron teletherapy
C0454077|T061|Teleradiotherapy using electrons
C0454077|T061|Electron teletherapy
C0278777|T061|Low-LET Cobalt-60 Gamma Ray Therapy
C1275217|T191|Paget Disease of the Vulva
C1275217|T191|Paget's Disease of Vulva
C1275217|T191|Vulvar Paget's Disease
C1275217|T191|Vulva Paget's Disease
C1275217|T191|Paget's Disease of the Vulva
CL378255|T061|Breathing-Synchronized Delivery Tomotherapy
CL378255|T061|BSD Tomotherapy
C1335759|T033|Resected Mass
C1335759|T033|Resectable Mass
C114761|T061|Intensity-Modulated Spot-Scanning Proton Therapy
C114761|T061|Spot Scan Intensity-Modulated Proton Therapy
C1300989|T201|Tumor size, largest metastasis
C1300989|T201|Tumour size, largest metastasis
C1300989|T201|Tumor size, largest metastasis (observable entity)
C0854810|T191|Recurrent Lymphocyte Depleted Classical Hodgkin Lymphoma
C0854810|T191|Relapsed Hodgkin's Disease Lymphocyte Depletion Type
C0854810|T191|Recurrent Hodgkin's Lymphoma Lymphocyte Depleted
C0854810|T191|Relapsed Hodgkin's Lymphoma Lymphocyte Depletion Type
C0854810|T191|Recurrent Hodgkin's Lymphoma Lymphocyte Depletion Type
C0854810|T191|Recurrent Hodgkin's Disease Lymphocyte Depletion Type
C0854810|T191|Hodgkin's disease lymphocyte depletion type recurrent
C0854810|T191|Recurrent Lymphocyte Depleted Hodgkin's Lymphoma
C0854810|T191|Recurrent Lymphocyte Depleted Hodgkin Lymphoma
C1333418|T191|Epipodophyllotoxin-Related Myelodysplastic Syndrome
C1333418|T191|Epipodophyllotoxin Related Myelodysplastic Syndrome
C1332261|T191|Paget Disease of the Anal Canal
C1332261|T191|Anal Canal Paget's Disease
C1332261|T191|Paget's Disease of the Anal Canal
C1332261|T191|Paget's Disease of Anal Canal
C0853971|T191|Stage IIIB Inflammatory Breast Carcinoma
C0853971|T191|Inflammatory Carcinoma of Breast Stage III
C0853971|T191|Stage III Inflammatory Breast Cancer
C0853971|T191|Stage III Inflammatory Breast Carcinoma
C0853971|T191|Stage IIIB Inflammatory Breast Cancer
C1708230|T033|Generic Distant Metastasis TNM Finding
C0730456|T170|Tumor stage T1mic
C0730456|T170|Tumor stage T1mic (finding)
C0730456|T170|Tumour stage T1mic
C3272501|T033|Ta Stage Finding
C0240225|T033|Hepatic Mass
C0240225|T033|LIVER MASS
C0240225|T033|Liver mass
C0240225|T033|mass
C0240225|T033|Liver Mass
C0240225|T033|Liver mass (finding)
C0240225|T033|liver mass
C0240225|T033|Hepatic mass
C1333008|T191|Childhood Testicular Mixed Embryonal Carcinoma and Teratoma
C1333008|T191|Childhood Teratocarcinoma of Testis
C1333008|T191|Childhood Testicular Teratocarcinoma
C1333008|T191|Pediatric Testicular Teratocarcinoma
C1333008|T191|Childhood Teratocarcinoma of the Testis
CL454083|T191|Classical Glioblastoma
C3272364|T033|T1mi Stage Finding
C0475372|T033|T1 Stage Finding
C0475372|T033|T1 Tumor Stage
C0475372|T033|T1 stage
C0475372|T033|Tumour stage T1
C0475372|T033|T1 TNM Finding
C0475372|T033|Tumor Stage T1
C0475372|T033|T1 Primary Tumor Finding
C0475372|T033|T1 category (finding)
C0475372|T033|Tumor stage T1
C0475372|T033|T1 category
C0475372|T033|T1
C0475372|T033|T1 Primary Tumor Stage Finding
C0475372|T033|T1 Tumor Finding
C0475372|T033|T1 Cancer Stage Finding
C0475372|T033|T1 tumor stage
C0475372|T033|T1 Stage
C0854744|T191|Stage I AIDS-Related Anal Canal Cancer
C0854744|T191|Stage I AIDS-Related Anal Canal Cancer AJCC v6
C0854744|T191|Stage I AIDS-Related Anal Canal Cancer AJCC v7
C3272458|T033|cM0 (i+) Stage Finding
C535972|T191|Lynch 1 Syndrome
C535972|T191|Syndrome, Lynch
C535972|T191|HNPCC - hereditary nonpolyposis colon cancer
C535972|T191|COLORECTAL CANCER, HEREDITARY NONPOLYPOSIS, TYPE 1
C535972|T191|Hereditary nonpolyposis colon cancer
C535972|T191|COCA1
C535972|T191|COLON CANCER, FAMILIAL NONPOLYPOSIS, TYPE 1
C535972|T191|Familial Non-Polyposis Colon Cancer Type 1
C535972|T191|HNPCC1
C535972|T191|Colon Cancer, Familial Nonpolyposis
C535972|T191|Colorectal Cancer Hereditary Nonpolyposis
C535972|T191|Colon cancer, familial nonpolyposis, type 1
C535972|T191|Hereditary Nonpolyposis Colorectal Cancer
C535972|T191|HNPCC
C535972|T191|Lynch Cancer Family Syndrome I
C535972|T191|FCC1
C535972|T191|Hereditary nonpolyposis colon cancer (disorder)
C535972|T191|Lynch Syndrome I
C535972|T191|Hereditary Nonpolyposis Colon Cancer
C535972|T191|LYNCH SYNDROME I
C535972|T191|Lynch Syndrome
C535972|T191|Colorectal cancer, hereditary nonpolyposis, type 1
C535972|T191|Hereditary Non-Polyposis Colon Cancer Type 1
C1335689|T191|Rectal Sarcomatoid Carcinoma
C1335689|T191|Rectal Spindle Cell Carcinoma
C1335689|T191|Sarcomatoid Carcinoma of the Rectum
C1335689|T191|Sarcomatoid Carcinoma of Rectum
C115093|T191|Recurrent Oropharyngeal Undifferentiated Carcinoma
C115093|T191|Oropharyngeal lymphoepithelioma recurrent
C115093|T191|lymphoepithelioma of the oropharynx, recurrent
C115093|T191|oropharyngeal lymphoepithelioma, recurrent
C115093|T191|recurrent lymphoepithelioma of the oropharynx
C115093|T191|Recurrent Oropharyngeal Lymphoepithelioma
C115093|T191|Oropharyngeal lymphepithelioma recurrent
C115093|T191|oropharynx lymphoepithelioma, recurrent
C0577691|T191|Disseminated Squamous Cell Carcinoma
C0577691|T191|Disseminated squamous cell carcinoma
C0577691|T191|Disseminated squamous cell carcinoma (morphologic abnormality)
C1333834|T191|Grade 1 Malignant Neoplasm
C1367874|T191|Metastatic Neoplasm of the Urethra
C1367874|T191|Metastatic Neoplasm of Urethra
C1367874|T191|Urethra Metastatic Malignant Neoplasm
C0877355|T191|Localized Gallbladder Carcinoma
C0877355|T191|Gallbladder Cancer, Localized
C0877355|T191|localized gallbladder cancer
C0877355|T191|Gallbladder carcinoma localized
C0877355|T191|Localized Gallbladder Cancer
C0877355|T191|gallbladder cancer, localized
C0877355|T191|Localized Cancer of the Gallbladder
C0877355|T191|Localized Cancer of Gallbladder
C0877355|T191|Gallbladder carcinoma localised
C0240318|T047|Mediastinal Mass
C0240318|T047|Mass of mediastinum (finding)
C0240318|T047|Mass of mediastinum
C0240318|T047|MEDIASTINAL MASS
C0240318|T047|Mediastinal mass
C0276535|T191|AIDS-Related Kaposi Sarcoma
C0276535|T191|Kaposi's Sarcoma Epidemic Type
C0276535|T191|Kaposi's Sarcoma AIDS Related
C0276535|T191|Autoimmune Deficiency Syndrome-Related Kaposi Sarcoma
C0276535|T191|AIDS-related Kaposi sarcoma
C0276535|T191|Epidemic Kaposi's Sarcoma
C0276535|T191|AIDS, Kaposi's Sarcoma
C0276535|T191|AIDS Related Kaposi's Sarcoma
C0276535|T191|AIDS-Related Kaposi's Sarcoma
C1334017|T191|High Grade Malignant Neoplasm
C0279017|T061|High-LET Heavy Ion Therapy
C0279017|T061|Therapy, High-LET Heavy Ion
C0279017|T061|Heavy Ion Radiation
C1301362|T191|Primary Cutaneous Anaplastic Large Cell Lymphoma
C1301362|T191|Anaplastic large-cell lymphoma, primary cutaneous type
C1301362|T191|Primary cutaneous CD30+ large T-cell lymphoma
C1301362|T191|Lymphoma, Primary Cutaneous Anaplastic Large Cell [Disease/Finding]
C1301362|T191|Primary cutaneous anaplastic large cell lymphoma
C1301362|T191|Primary cutaneous anaplastic large T-cell lymphoma, CD30-positive (morphologic abnormality)
C1301362|T191|Cutaneous T-cell lymphoma, large cell, CD30-positive
C1301362|T191|Primary cutaneous CD30 antigen positive large T-cell lymphoma (disorder)
C1301362|T191|Primary cutaneous CD30-positive large T-cell lymphoma
C1301362|T191|ALCL, cutaneous
C1301362|T191|Primary Anaplastic Large Cell Lymphoma of the Skin
C1301362|T191|Primary Cutaneous CD30+ Anaplastic Large Cell Lymphoma
C1301362|T191|Primary Cutaneous CD30 positive Large T Cell Lymphoma
C1301362|T191|Lymphoma, Primary Cutaneous Anaplastic Large Cell
C1301362|T191|Primary Cutaneous CD30 Positive Anaplastic Large Cell Lymphoma
C1301362|T191|Primary Cutaneous CD30+ ALCL
C1301362|T191|C-ALCL
C1301362|T191|Primary cutaneous anaplastic large T-cell lymphoma, CD30-positive
C1301362|T191|Anaplastic large-cell lymphoma, primary cutaneous type 
C1301362|T191|Anaplastic large cell lymphoma, T/Null cell, primary cutaneous type
C1301362|T191|Primary Anaplastic Large Cell Lymphoma of Skin
C1301362|T191|Primary cutaneous CD30 antigen positive large T-cell lymphoma
C1301362|T191|Anaplastic large cell lymphoma, cutaneous type
C1301362|T191|Primary Cutaneous CD30-positive Large T-Cell Lymphoma
C1301362|T191|Primary cutaneous CD30-positive T-cell proliferations
CL433949|T191|Recurrent Childhood Anaplastic Oligoastrocytoma
CL433949|T191|recurrent childhood anaplastic oligoastrocytoma
C0278519|T191|Recurrent Childhood Acute Lymphoblastic Leukemia
C0278519|T191|Recurrent Pediatric Acute Lymphocytic Leukemia
C0278519|T191|recurrent childhood ALL
C0278519|T191|ALL, recurrent, childhood
C0278519|T191|Relapsed Pediatric Acute Lymphocytic Leukemia
C0278519|T191|Recurrent Pediatric ALL
C0278519|T191|childhood ALL, recurrent
C0278519|T191|recurrent childhood acute lymphoblastic leukemia
C0278519|T191|relapsed pediatric acute lymphocytic leukemia
C0278519|T191|relapsed pediatric ALL
C0278519|T191|Recurrent Pediatric Acute Lymphoid Leukemia
C0278519|T191|Relapsed Pediatric ALL
C0278519|T191|Recurrent Childhood Acute Lymphocytic Leukemia
C0278519|T191|recurrent pediatric acute lymphogenous leukemia
C0278519|T191|Relapsed Childhood ALL
C0278519|T191|Relapsed Pediatric Acute Lymphogenous Leukemia
C0278519|T191|recurrent childhood acute lymphoid leukemia
C0278519|T191|Recurrent Childhood Precursor Lymphoblastic Leukemia
C0278519|T191|acute lymphocytic leukemia, childhood, relapsed
C0278519|T191|Relapsed Childhood Acute Lymphoblastic Leukemia
C0278519|T191|Relapsed Pediatric Acute Lymphoid Leukemia
C0278519|T191|recurrent childhood acute lymphogenous leukemia
C0278519|T191|ALL, recurrent, pediatric
C0278519|T191|ALL, pediatric, relapsed
C0278519|T191|relapsed childhood acute lymphoblastic leukemia
C0278519|T191|Relapsed Childhood Acute Lymphocytic Leukemia
C0278519|T191|relapsed childhood ALL
C0278519|T191|recurrent pediatric ALL
C0278519|T191|childhood acute lymphocytic leukemia, relapsed
C0278519|T191|ALL, relapsed, pediatric
C0278519|T191|pediatric acute lymphocytic leukemia, relapsed
C0278519|T191|relapsed pediatric acute lymphoblastic leukemia
C0278519|T191|Relapsed Pediatric Acute Lymphoblastic Leukemia
C0278519|T191|relapsed childhood acute lymphocytic leukemia
C0278519|T191|Recurrent Childhood ALL
C0278519|T191|lymphocytic leukemia, acute, childhood, relapsed
C0278519|T191|childhood ALL, relapsed
C0278519|T191|relapsed pediatric acute lymphogenous leukemia
C0278519|T191|relapsed pediatric acute lymphoid leukemia
C0278519|T191|ALL, relapsed, childhood
C0278519|T191|Recurrent Pediatric Acute Lymphoblastic Leukemia
C0278519|T191|recurrent pediatric acute lymphocytic leukemia
C0278519|T191|Recurrent Pediatric Acute Lymphogenous Leukemia
C0278519|T191|leukemia, acute lymphocytic, childhood, relapsed
C0278519|T191|pediatric ALL, recurrent
C0278519|T191|pediatric ALL, relapsed
C0278519|T191|Recurrent Childhood Acute Lymphoid Leukemia
C0278519|T191|ALL, childhood, relapsed
C0278519|T191|recurrent pediatric acute lymphoblastic leukemia
C0278519|T191|recurrent childhood precursor lymphoblastic leukemia
C0278519|T191|recurrent pediatric acute lymphoid leukemia
C0278519|T191|Recurrent Childhood Acute Lymphogenous Leukemia
C0279028|T061|Ablative Endocrine Surgery
C0279028|T061|ablative endocrine surgery
C0279028|T061|surgery, ablative endocrine
CL472796|T191|Recurrent Malignant Extragonadal Germ Cell Tumor
C0279986|T191|Childhood Leiomyosarcoma
C0279986|T191|leiomyosarcoma, childhood
C0279986|T191|sarcoma, leiomyo-, childhood
C0279986|T191|sarcoma, leiomyo-, pediatric
C0279986|T191|Pediatric Leiomyosarcoma
C0279986|T191|leiomyosarcoma, pediatric
C0279986|T191|pediatric leiomyosarcoma
C0279986|T191|childhood leiomyosarcoma
C1335513|T191|Acinar Prostate Mucinous Adenocarcinoma
C1335513|T191|Colloidal Prostate Adenocarcinoma
C1335513|T191|Colloidal Adenocarcinoma of the Prostate
C1335513|T191|Colloidal Adenocarcinoma of Prostate
C1335513|T191|Colloid Adenocarcinoma of the Prostate
C1335513|T191|Acinar Colloid Prostate Adenocarcinoma
C1335513|T191|Colloid Adenocarcinoma of Prostate
C1335513|T191|Mucinous Adenocarcinoma of the Prostate
C1335513|T191|Mucinous Adenocarcinoma of Prostate
C0347012|T191|Metastatic Malignant Neoplasm to the Urethra
C0347012|T191|Metastasis to the Urethra
C0347012|T191|Metastatic Neoplasm to the Urethra
C120286|T081|Tumor Greater Than or Equal to 2.1 Centimeters
C120286|T081|Greater than or equal to 2.1 cm
C1332898|T191|Centroblastic Lymphoma Post-Transplant Lymphoproliferative Disorder
C1332898|T191|Centroblastic Lymphoma PTLD
C1332898|T191|Centroblastic Diffuse Large B-Cell Lymphoma PTLD
C0442835|T046|Atypical Lobular Breast Hyperplasia
C0442835|T046|Atypical Lobular Hyperplasia of Breast
C0442835|T046|atypical lobular hyperplasia of the breast
C0442835|T046|atypical lobular hyperplasia
C0442835|T046|Atypical lobular hyperplasia of breast (disorder)
C0442835|T046|atypical breast lobular hyperplasia
C0442835|T046|Atypical Lobular Hyperplasia of the Breast
C0442835|T046|atypical lobular hyperplasia of breast
C0442835|T046|Atypical lobular hyperplasia of breast
C0442835|T046|ALH
C0442835|T046|Atypical Breast Lobular Hyperplasia
C0442835|T046|atypical lobular breast hyperplasia
C0442835|T046|Atypical lobular hyperplasia
C0442835|T046|Atypical lobular hyperplasia (morphologic abnormality)
C1321869|T191|Childhood Intraocular Retinoblastoma
C1321869|T191|pediatric intraocular retinoblastoma
C1321869|T191|childhood intraocular retinoblastoma
C1321869|T191|Pediatric Intraocular Retinoblastoma
C0854970|T191|Recurrent Adenosquamous Lung Carcinoma
C0854970|T191|Adenosquamous Cell Lung Carcinoma Recurrent
C0854970|T191|Adenosquamous cell lung cancer recurrent
C0854970|T191|Recurrent Adenosquamous Cell Lung Carcinoma
C0854970|T191|Recurrent Adenosquamous Cell Carcinoma of the Lung
C0854970|T191|Recurrent Adenosquamous Cell Carcinoma of Lung
C1541449|T191|Recurrent Grade II Lymphomatoid Granulomatosis
C1880431|T061|E-CMF Regimen
C1880431|T061|Epirubicin-Cytoxan-Methotrexate-Fluorouracil Regimen
C0587052|T033|Hilar Mass
C0587052|T033|Pulmonary Hilum Mass
C0587052|T033|Mass of hilum
C0587052|T033|Pulmonary hilum mass
C0587052|T033|Hilar mass
C0587052|T033|Mass of hilum (finding)
C1709110|T033|N3c Stage Finding
C1709110|T033|N3c Cancer Stage Finding
C1709110|T033|N3c Node Finding
C1709110|T033|N3c Lymph Node Stage
C1709110|T033|N3c Node Stage
C1709110|T033|N3c Lymph Node Finding
C1709110|T033|N3c
C1709110|T033|N3c Regional Lymph Nodes Finding
C1709110|T033|N3c Regional Lymph Node Stage Finding
C1709110|T033|N3c TNM Finding
C1709110|T033|Node Stage N3c
C1709110|T033|N3c Stage
C1709110|T033|Lymph Node Stage N3c
C1881358|T033|Large Mass
C1519370|T191|Anaplastic Large Cell Lymphoma, Signet Ring-Like Subtype
C0854178|T191|Metastatic Malignant Neoplasm to the Adrenal Gland
C0854178|T191|Metastatic Tumor to the Adrenals
C0854178|T191|Metastasis to Adrenals
C0854178|T191|Metastatic Neoplasm to the Adrenal Gland
C0854178|T191|Metastatic Tumor to the Adrenal Gland
C0854178|T191|Metastases to Adrenals
C0854178|T191|Metastatic Neoplasm to the Adrenals
C0751623|T191|Secondary Malignant Neoplasm
C0751623|T191|Second Primary Cancer
C0751623|T191|Treatment related secondary malignancy
C0751623|T191|Secondary Cancer
C0751623|T191|Cancer, Second
C0751623|T191|secondary cancer
C0751623|T191|Second Primary Cancers
C0751623|T191|Second Cancers
C0751623|T191|Cancer, Second Primary
C0751623|T191|Cancers, Second Primary
C0751623|T191|Secondary Malignancy
C0751623|T191|Second Cancer
C0751623|T191|Cancers, Second
C0751623|T191|Second primary malignancy
C1515862|T191|Acinar Prostate Adenocarcinoma, Atrophic Variant
C0280788|T191|Anaplastic Ependymoma
C0280788|T191|anaplastic ependymoma (WHO grade III)
C0280788|T191|anaplastic ependymoma
C0280788|T191|EPENDYMOMA, ANAPLASTIC , MALIGNANT
C0280788|T191|Ependymoma, anaplastic (morphologic abnormality)
C0280788|T191|Anaplastic ependymoma
C0280788|T191|ANAPLASTIC EPENDYMAL NEOPLASM
C0280788|T191|Malignant Ependymoma
C0280788|T191|WHO Grade III Ependymal Tumor
C0280788|T191|MALIGNANT EPENDYMOMA
C0280788|T191|Anaplastic Ependymal Neoplasm
C0280788|T191|UNDIFFERENTIATED EPENDYMOMA
C0280788|T191|Undifferentiated Ependymal Tumor
C0280788|T191|UNDIFFERENTIATED EPENDYMAL NEOPLASM
C0280788|T191|Ependymomas, Anaplastic
C0280788|T191|Ependymoma, anaplastic
C0280788|T191|Ependymoma malignant
C0280788|T191|WHO Grade III Ependymal Neoplasm
C0280788|T191|Anaplastic Ependymomas
C0280788|T191|ependymoma (WHO grade III)
C0280788|T191|UNDIFFERENTIATED EPENDYMAL TUMOR
C0280788|T191|WHO GRADE III EPENDYMAL TUMOR
C0280788|T191|ANAPLASTIC EPENDYMAL TUMOR
C0280788|T191|WHO GRADE III EPENDYMAL NEOPLASM
C0280788|T191|Anaplastic Ependymal Tumor
C0280788|T191|Undifferentiated Ependymoma
C0280788|T191|Undifferentiated Ependymal Neoplasm
C0280788|T191|Ependymoma, Anaplastic
C1705427|T045|Germline Mutation
C1705427|T045|Germline Mutations
C1705427|T045|Mutation, Germline
C1705427|T045|Germ Line Mutation
C1705427|T045|Mutation, Germ-Line
C1705427|T045|germline mutation
C1705427|T045|Mutations, Germline
C1705427|T045|Mutations, Germ-Line
C1705427|T045|Hereditary Mutation
C1705427|T045|Germ-Line Mutation
C1705427|T045|hereditary mutation
C1705427|T045|Germline Mutation Abnormality
C1705427|T045|Germ-Line Mutations
C1705427|T045|Mutation, Germ Line
C0278704|T191|Malignant Childhood Neoplasm
C0278704|T191|pediatric cancer
C0278704|T191|Malignant Pediatric Tumor
C0278704|T191|childhood cancer
C0278704|T191|pediatric neoplasm
C0278704|T191|Malignant Pediatric Neoplasm
C0278704|T191|Malignant Childhood Tumor
C0278704|T191|Pediatric Cancer
C0278704|T191|cancer, childhood
C0278704|T191|Childhood Cancer
C0278704|T191|pediatric neoplasm/cancer
CL378277|T061|Humidification-Modulated Radiation Therapy
C0686463|T191|Metastatic Malignant Neoplasm to the Ciliary Body
C0686463|T191|Metastatic Neoplasm to the Ciliary Body
C0686463|T191|Metastatic Tumor to the Ciliary Body
C0686463|T191|Metastasis to the Ciliary Body
C0279566|T191|Paget Disease and Intraductal Carcinoma of the Breast
C0279566|T191|Paget's Disease of the Breast with Intraductal Carcinoma
C0279566|T191|Paget's Disease of Breast with Intraductal Carcinoma
C0279566|T191|Paget's Disease and Intraductal Carcinoma of the Breast
C0279566|T191|Paget's Disease and Intraductal Carcinoma of Breast
C0600521|T061|3-Dimensional Conformal Radiation Therapy
C0600521|T061|Radiation Conformal Therapy
C0600521|T061|3-dimensional radiation therapy
C0600521|T061|3D-CRT
C0600521|T061|Conformal Therapy
C0600521|T061|3-dimensional conformal radiation therapy
C1335476|T191|Central Nervous System Anaplastic Large Cell Lymphoma
C1335476|T191|Anaplastic Large Cell Lymphoma of Central Nervous System
C1335476|T191|Anaplastic Central Nervous System Large Cell Lymphoma
C1335476|T191|Primary Central Nervous System Anaplastic Large Cell Lymphoma
C1335476|T191|Anaplastic Large Cell Lymphoma of CNS
C1335476|T191|Anaplastic Large Cell Lymphoma of the CNS
C1335476|T191|Anaplastic CNS Large Cell Lymphoma
C1335476|T191|Anaplastic Large Cell Lymphoma of the Central Nervous System
C1335476|T191|Primary CNS Anaplastic Large Cell Lymphoma
C0278779|T191|Recurrent Osteosarcoma
C0278779|T191|recurrent osteosarcoma
C0278779|T191|recurrent osteogenic sarcoma
C0278779|T191|Osteosarcoma recurrent
C0278779|T191|osteogenic sarcoma, recurrent
C0278779|T191|sarcoma, recurrent osteogenic
C0278779|T191|Osteogenic sarcoma recurrent
C0278779|T191|Relapsed Osteogenic Sarcoma
C0278779|T191|osteosarcoma, recurrent
C0278779|T191|Recurrent Osteogenic Sarcoma
C0278779|T191|Osteosarcoma, Recurrent
C0278779|T191|Relapsed Osteosarcoma
C116430|T061|4-Dimensional Conformal Radiation Therapy
C116430|T061|4D Conformal Radiation Therapy
C0203608|T061|Isotope Therapy
C0203608|T061|radionuclide therapy
C0203608|T061|Radionuclide therapy
C0203608|T061|Radionuclide therapy (procedure)
C0203608|T061|Radioactive Isotope Therapy
C0203608|T061|Internal radiotherapy
C0203608|T061|Radioisotope Therapy
C0203608|T061|Radioisotope therapy
C0203608|T061|Short distance and contact radiotherapy
C0203608|T061|RI - Radioisotope therapy
C0203608|T061|radioactive isotope therapy
C0203608|T061|radioisotope therapy
C0203608|T061|Radiotherapy - internal
C0203608|T061|therapy, isotope, radioactive
C0203608|T061|Radioisotope teleradiotherapy
C0278698|T191|Stage III Childhood Hepatocellular Carcinoma
C0278698|T191|Stage III Pediatric Hepatoma
C0278698|T191|Stage III Childhood Hepatoma
C0278698|T191|Stage III Pediatric Liver Cell Carcinoma
C0278698|T191|Stage III Childhood Hepatocellular Carcinoma AJCC v7
C0278698|T191|Stage III Pediatric Hepatocellular Carcinoma
C0278698|T191|Stage III Childhood Liver Cell Carcinoma
C0278698|T191|stage III childhood liver cancer
C0279918|T191|Recurrent Childhood Hodgkin Lymphoma
C0279918|T191|relapsed Hodgkin's disease, childhood
C0279918|T191|HD, pediatric, recurrent
C0279918|T191|Recurrent Childhood Hodgkin's Disease
C0279918|T191|childhood HD, recurrent
C0279918|T191|HD, childhood, relapsed
C0279918|T191|childhood HD, relapsed
C0279918|T191|recurrent HD, pediatric
C0279918|T191|pediatric Hodgkin's disease, relapsed
C0279918|T191|Hodgkin's lymphoma, relapsed, childhood
C0279918|T191|relapsed pediatric Hodgkin's disease
C0279918|T191|recurrent HD, childhood
C0279918|T191|Relapsed Childhood Hodgkin's Disease
C0279918|T191|Recurrent Pediatric Hodgkin's Disease
C0279918|T191|HD, childhood, recurrent
C0279918|T191|recurrent pediatric HD
C0279918|T191|Hodgkin's disease, recurrent, childhood
C0279918|T191|recurrent childhood HD
C0279918|T191|Relapsed Childhood Hodgkin's Lymphoma
C0279918|T191|lymphoma, relapsed childhood Hodgkin's
C0279918|T191|refractory childhood Hodgkin's disease
C0279918|T191|relapsed HD, childhood
C0279918|T191|childhood Hodgkin's disease, relapsed
C0279918|T191|recurrent/refractory childhood Hodgkin lymphoma
C0279918|T191|relapsed childhood Hodgkin's disease
C0279918|T191|relapsed childhood HD
C0279918|T191|Recurrent Pediatric Hodgkin's Lymphoma
C0279918|T191|HD, childhood, refractory
C0279918|T191|refractory childhood HD
C0279918|T191|recurrent/refractory childhood Hodgkin's disease
C0279918|T191|HD, relapsed, childhood
C0279918|T191|Hodgkin's disease, relapsed, childhood
C0279918|T191|Relapsed Pediatric Hodgkin's Disease
C0279918|T191|pediatric HD, relapsed
C0279918|T191|recurrent pediatric Hodgkin's disease
C0279918|T191|Recurrent Childhood Hodgkin's Lymphoma
C0279918|T191|Relapsed Pediatric Hodgkin's Lymphoma
C0279918|T191|recurrent Hodgkin's disease, childhood
C1711365|T061|Limited Radiation Therapy
C0475390|T185|T3a Stage Finding
C0475390|T185|Tumor stage T3a
C0475390|T185|Tumor stage T3a (finding)
C0475390|T185|Tumour stage T3a
C0475390|T185|T3a Cancer Stage Finding
C0475390|T185|T3a TNM Finding
C0475390|T185|T3a tumor stage
C0475390|T185|T3a Primary Tumor Stage Finding
C0475390|T185|T3a
C0475390|T185|T3a Tumor Finding
C0475390|T185|T3a Stage
C0475390|T185|T3a Tumor Stage
C0475390|T185|T3a Primary Tumor Finding
C0475390|T185|Tumor Stage T3a
C0278778|T061|Low-LET Photon Therapy
C1541448|T191|Recurrent Grade I Lymphomatoid Granulomatosis
C0279583|T191|Childhood T Acute Lymphoblastic Leukemia
C0279583|T191|T-Cell Childhood Acute Lymphoblastic Leukemia
C0279583|T191|T-Cell Childhood ALL
C0279583|T191|T-Cell Pediatric Acute Lymphocytic Leukemia
C0279583|T191|T-Cell Pediatric Acute Lymphoblastic Leukemia
C0279583|T191|Childhood Precursor T-Lymphoblastic Leukemia
C0279583|T191|T-Cell Childhood Acute Lymphocytic Leukemia
C0279583|T191|T-Cell Pediatric ALL
C0279583|T191|Childhood T-Cell Acute Lymphoblastic Leukemia
C0347010|T191|Metastatic Malignant Neoplasm to the Ureter
C0347010|T191|Metastatic Neoplasm to the Ureter
C0347010|T191|Metastatic Tumor to the Ureter
C0347010|T191|Metastasis to the Ureter
C0206180|T191|Anaplastic Large Cell Lymphoma
C0206180|T191|LYMPHOMA LARGE CELL KI 01
C0206180|T191|CD 030 POSITIVE ANAPLASTIC LARGE CELL LYMPHOMA
C0206180|T191|Lymphoma, Large-Cell, Anaplastic [Disease/Finding]
C0206180|T191|Anaplastic large cell lymphoma T- and null-cell types
C0206180|T191|Systemic Anaplastic Large-Cell Lymphoma
C0206180|T191|Anaplastic large cell lymphoma, CD30-positive
C0206180|T191|Anaplastic large cell lymphoma, CD30+
C0206180|T191|Ki-1 Lymphoma
C0206180|T191|Anaplastic large cell lymphoma (ALCL) CD30+
C0206180|T191|anaplastic large cell lymphoma
C0206180|T191|Anaplastic large cell lymphoma, NOS
C0206180|T191|Systemic Anaplastic Large Cell Lymphoma
C0206180|T191|(Ki-1+) lymphoma
C0206180|T191|Large cell (Ki-1+) lymphoma [obs]
C0206180|T191|Anaplastic large cell lymphoma T- and null-cell types NOS
C0206180|T191|ANAPLASTIC LARGE CELL LYMPHOMA
C0206180|T191|Ki 1 Lymphoma
C0206180|T191|Large-Cell Lymphoma, Anaplastic
C0206180|T191|Ki-1+ ALCL
C0206180|T191|Anaplastic Large-Cell Lymphoma
C0206180|T191|CD30+ Anaplastic Large-Cell Lymphoma
C0206180|T191|Lymphoma, Large-Cell, Anaplastic
C0206180|T191|Lymphoma, Anaplastic Large-Cell
C0206180|T191|Large-Cell Lymphomas, Anaplastic
C0206180|T191|Ki-1 Lymphomas
C0206180|T191|Lymphomas, Ki-1
C0206180|T191|CD30 Positive Anaplastic Large Cell Lymphoma
C0206180|T191|lymphoma, anaplastic large cell
C0206180|T191|Lymphoma, Large-Cell, Ki-1
C0206180|T191|Anaplastic large cell lymphomas T- and null-cell types
C0206180|T191|Anaplastic Large-Cell Lymphomas
C0206180|T191|Anaplastic large cell lymphoma
C0206180|T191|Anaplastic large-cell lymphoma
C0206180|T191|Large cell anaplastic lymphoma (disorder)
C0206180|T191|Ki-1+ Anaplastic Large Cell Lymphoma
C0206180|T191|ALCL
C0206180|T191|CD30-Positive Anaplastic Large-Cell Lymphoma
C0206180|T191|Large cell anaplastic lymphoma
C0206180|T191|Lymphoma, Ki-1
C0206180|T191|CD30+ Anaplastic Large Cell Lymphoma
C0206180|T191|Lymphomas, Anaplastic Large-Cell
C0206180|T191|Anaplastic large cell lymphoma, T cell and Null cell type (morphologic abnormality)
C0206180|T191|Anaplastic large cell lymphoma, T cell and Null cell type
C1514511|T191|Prostate Ductal Adenocarcinoma, Cribriform Pattern
C0007344|T061|Surgical Castration
C0007344|T061|surgical castration
C0007344|T061|Castration
C0007344|T061|castration
C0007344|T061|CASTRATION
C0007344|T061|Castrations
C1334745|T191|Methotrexate-Associated Burkitt Lymphoma
C1334745|T191|Methotrexate-Associated Burkitt's Lymphoma
C1333981|T191|Hepatoblastoma with Combined Fetal and Embryonal Epithelial Differentiation
C0347011|T191|Metastatic Malignant Neoplasm to the Bladder
C0347011|T191|Metastatic Neoplasm to the Urinary Bladder
C0347011|T191|Metastases to Bladder
C0347011|T191|Metastatic Tumor to the Bladder
C0347011|T191|Metastatic Neoplasm to the Bladder
C0347011|T191|Metastasis to Bladder
C0347011|T191|Metastatic Tumor to the Urinary Bladder
C115429|T191|Recurrent Fallopian Tube Carcinoma
C0744049|T047|Flank Mass
C0804677|T082|Tumor size
C0804677|T082|tumor size
C0804677|T082|Tumor size (observable entity)
C0804677|T082|Size:Len:Pt:Tumor:Qn
C0804677|T082|Size Tumor
C0804677|T082|size of tumor
C0804677|T082|Size:Length:Point in time:Tumor:Quantitative
C0804677|T082|Tumour size
C0804677|T082|Size of tumor
C0804677|T082|Size of tumour
C0280449|T191|Secondary Acute Myeloid Leukemia
C0280449|T191|secondary AML
C0280449|T191|secondary acute non-lymphocytic leukemia
C0280449|T191|secondary acute nonlymphoblastic leukemia
C0280449|T191|Secondary AGL
C0280449|T191|Secondary Acute Myeloblastic Leukemia
C0280449|T191|Secondary Acute Granulocytic Leukemia
C0280449|T191|acute nonlymphocytic leukemia, secondary
C0280449|T191|nonlymphocytic leukemia, secondary acute
C0280449|T191|acute non-lymphoblastic leukemia, secondary
C0280449|T191|Secondary AML
C0280449|T191|Secondary Acute Myelocytic Leukemia
C0280449|T191|non-lymphoblastic leukemia, secondary acute
C0280449|T191|secondary acute non-lymphoblastic leukemia
C0280449|T191|acute nonlymphoblastic leukemia, secondary
C0280449|T191|acute non-lymphocytic leukemia, secondary
C0280449|T191|secondary acute myelogenous leukemia
C0280449|T191|secondary ANLL
C0280449|T191|nonlymphoblastic leukemia, secondary acute
C0280449|T191|acute myelogenous leukemia, secondary
C0280449|T191|myelogenous leukemia, secondary acute
C0280449|T191|secondary acute myeloid leukemia
C0280449|T191|non-lymphocytic leukemia, secondary acute
C0280449|T191|secondary acute nonlymphocytic leukemia
C0280449|T191|acute myeloid leukemia, secondary
C0280449|T191|Secondary Acute Myelogenous Leukemia
C0280449|T191|myeloid leukemia, secondary acute
C115966|T191|Infiltrating Bladder Urothelial Carcinoma Associated with Urethral Carcinoma
C0279987|T191|Childhood Malignant Peripheral Nerve Sheath Tumor
C0279987|T191|neurolemma, malignant, childhood
C0279987|T191|Childhood Malignant Neoplasm of Peripheral Nerve Sheath
C0279987|T191|Childhood Malignant Tumor of the Peripheral Nerve Sheath
C0279987|T191|Childhood MPNST
C0279987|T191|Pediatric Malignant Peripheral Nerve Sheath Tumor
C0279987|T191|neurogenic sarcoma, childhood
C0279987|T191|Pediatric Malignant Schwannoma
C0279987|T191|Childhood Malignant Schwannoma
C0279987|T191|Pediatric MPNST
C0279987|T191|Pediatric Malignant Neurilemmoma
C0279987|T191|Pediatric Malignant Neoplasm of Peripheral Nerve Sheath
C0279987|T191|childhood neurofibrosarcoma
C0279987|T191|Childhood Malignant Tumor of Peripheral Nerve Sheath
C0279987|T191|Pediatric Malignant Peripheral Nerve Sheath Neoplasm
C0279987|T191|Childhood Malignant Neoplasm of the Peripheral Nerve Sheath
C0279987|T191|sarcoma, neurogenic, childhood
C0279987|T191|Childhood Malignant Neurilemmoma
C0279987|T191|Pediatric Malignant Neoplasm of the Peripheral Nerve Sheath
C0279987|T191|schwannoma, malignant, childhood
C0279987|T191|pediatric neurofibrosarcoma
C0279987|T191|sarcoma, neurofibro-, childhood
C0279987|T191|Pediatric Malignant Tumor of Peripheral Nerve Sheath
C0279987|T191|malignant neurolemma, childhood
C0279987|T191|malignant schwannoma, childhood
C0279987|T191|neurofibrosarcoma, pediatric
C0279987|T191|Childhood Malignant Peripheral Nerve Sheath Neoplasm
C0279987|T191|Pediatric Malignant Tumor of the Peripheral Nerve Sheath
C0279987|T191|neurofibrosarcoma, childhood
C116435|T061|3-Dimensional Conformal Accelerated Partial Breast Irradiation
C116435|T061|3D Conformal Accelerated Partial Breast Irradiation
C0205699|T191|Carcinomatosis
C0205699|T191|CARCINOMATOSIS
C0205699|T191|Carcinomatoses
C0205699|T191|carcinomatosis
C0205699|T191|Disseminated carcinomatosis
C0205699|T191|Carcinomatosis (morphologic abnormality)
C0205699|T191|Carcinomatosis (disorder)
C0205699|T191|carcinosis
C0205699|T191|[M]Carcinomatosis
C0205699|T191|Carcinomatosis NOS
C0677723|T191|Recurrent Indolent Adult Non-Hodgkin Lymphoma
C0677723|T191|Recurrent Adult Indolent Non-Hodgkin's Lymphoma
C0677723|T191|Recurrent Indolent Adult Non-Hodgkin's Lymphoma
CL383485|T191|Childhood Ependymoblastoma
CL383485|T191|childhood ependymoblastoma
CL433918|T191|Recurrent Childhood Gliosarcoma
CL433918|T191|recurrent childhood gliosarcoma
C1332625|T191|Breast Carcinoma Metastatic to the Liver
C1333293|T191|Diffuse Large B-Cell Lymphoma Post-Transplant Lymphoproliferative Disorder
C1333293|T191|Diffuse Large B-Cell Lymphoma PTLD
CL378646|T061|Total Marrow Irradiation
CL378646|T061|TMI
CL378646|T061|total marrow irradiation
C1299215|T201|Polyp size, dimension 3
C1299215|T201|Polyp size, dimension 3 (observable entity)
C1710405|T049|Thymidine to Cytosine Transition Abnormality
C1710405|T049|Thymidine to Cytosine Mutation
C1710405|T049|Thymidine to Cytosine Transition
C0036132|T061|Salpingo-Oophorectomy
C0036132|T061|salpingo-oophorectomy
C0854964|T191|Recurrent Penile Carcinoma
C0854964|T191|Relapsed Carcinoma of Penis
C0854964|T191|Penis carcinoma recurrent
C0854964|T191|Recurrent Penis Cancer
C0854964|T191|Recurrent Penile Cancer
C0854964|T191|Recurrent Penis Carcinoma
C0854964|T191|Relapsed Carcinoma of the Penis
C0854964|T191|recurrent penile cancer
C0854964|T191|penis cancer, recurrent
C0854964|T191|Relapsed Penile Carcinoma
C0854964|T191|Recurrent Carcinoma of Penis
C0854964|T191|Recurrent Carcinoma of the Penis
C0854964|T191|penile cancer, recurrent
C1336925|T191|AIDS-Related Gastric Kaposi Sarcoma
C1336925|T191|AIDS-Related Kaposi's Sarcoma of the Stomach
C1336925|T191|AIDS-Related Gastric Kaposi's Sarcoma
C1336925|T191|AIDS-Related Kaposi's Sarcoma of Stomach
C1299213|T201|Polyp size, dimension 1
C1299213|T201|Polyp size, dimension 1 (observable entity)
C1299214|T201|Polyp size, dimension 2
C1299214|T201|Polyp size, dimension 2 (observable entity)
C0281267|T191|Bilateral Breast Carcinoma
C0281267|T191|bilateral breast cancer
C0281267|T191|bilateral
C0281267|T191|Bilateral Breast Cancer
C0279615|T191|Childhood Mixed Alveolar Rhabdomyosarcoma
C0279615|T191|Pediatric Mixed Rhabdomyosarcoma
C0279615|T191|mixed cell type childhood rhabdomyosarcoma
C0279615|T191|Pediatric Mixed Type Rhabdomyosarcoma
C0279615|T191|rhabdomyosarcoma, mixed childhood
C0279615|T191|childhood rhabdomyosarcoma, mixed
C0279615|T191|rhabdomyosarcoma, pediatric mixed
C0279615|T191|mixed type pediatric rhabdomyosarcoma
C0279615|T191|pediatric rhabdomyosarcoma, mixed
C0279615|T191|rhabdomyosarcoma, childhood mixed
C0279615|T191|Childhood Mixed Cell Type Rhabdomyosarcoma
C0279615|T191|mixed cell type pediatric rhabdomyosarcoma
C0279615|T191|Childhood Mixed Type Rhabdomyosarcoma
C0279615|T191|mixed childhood rhabdomyosarcoma
C0279615|T191|Mixed Childhood Rhabdomyosarcoma
C0279615|T191|mixed pediatric rhabdomyosarcoma
C0279615|T191|Pediatric Mixed Cell Type Rhabdomyosarcoma
C0279615|T191|mixed type childhood rhabdomyosarcoma
C0280185|T191|Recurrent Grade 3 Follicular Lymphoma
C0280185|T191|follicular large cell lymphoma, relapsed
C0280185|T191|Relapsed Follicular Large Cell Lymphoma
C0280185|T191|Recurrent Grade III Follicular Large Cell Lymphoma
C0280185|T191|relapsed follicular large cell lymphoma
C0280185|T191|Relapsed Grade III Follicular Lymphoma
C0280185|T191|Recurrent Grade III Follicular Lymphoma
C0280185|T191|follicular large cell lymphoma, recurrent
C0280185|T191|recurrent grade 3 follicular lymphoma
C0280185|T191|Recurrent Follicular Large Cell Lymphoma
C0280185|T191|Relapsed Grade III Follicular Large Cell Lymphoma
C0280185|T191|recurrent grade III follicular large cell lymphoma
C1332642|T191|Burkitt-Like Lymphoma Post-Transplant Lymphoproliferative Disorder
C1332642|T191|Burkitt's-Like Lymphoma Post-Transplant Lymphoproliferative Disorder
C1332642|T191|Burkitt's-like Lymphoma PTLD
C1332642|T191|Burkitt-like Lymphoma PTLD
C1832047|T061|Balloon Brachytherapy
C1832047|T061|balloon catheter radiation
C1832047|T061|MammoSite
C0855012|T191|Metastatic Chondrosarcoma
C0855012|T191|Chondrosarcoma metastatic
C0855012|T191|Chondrosarcoma, Metastatic
C0279921|T191|Childhood Nodular Sclerosis Classical Hodgkin Lymphoma
C0279921|T191|Pediatric Nodular Sclerosis Hodgkin's Disease
C0279921|T191|pediatric nodular sclerosis Hodgkin's disease
C0279921|T191|childhood Hodgkin's disease, nodular sclerosis
C0279921|T191|Childhood NSHD
C0279921|T191|Pediatric Hodgkin's Nodular Sclerosis
C0279921|T191|Hodgkin's disease, nodular sclerosis, childhood
C0279921|T191|Childhood Hodgkin's Nodular Sclerosis
C0279921|T191|Childhood Nodular Sclerosis Hodgkin Lymphoma
C0279921|T191|pediatric HD, nodular sclerosis
C0279921|T191|Childhood Nodular Sclerosis Hodgkin's Lymphoma
C0279921|T191|Pediatric NSHD
C0279921|T191|Childhood Nodular Sclerosis Hodgkin's Disease
C0279921|T191|nodular sclerosing HD, childhood
C0279921|T191|nodular sclerosis Hodgkin's disease, childhood
C0279921|T191|pediatric Hogkin's disease, nodular sclerosis
C0279921|T191|Pediatric Nodular Sclerosis Hodgkin's Lymphoma
C0279921|T191|childhood nodular sclerosis Hodgkin's disease
C0279921|T191|childhood HD, nodular sclerosis
C0279921|T191|childhood nodular sclerosis Hodgkin lymphoma
C0279921|T191|nodular sclerosing Hodgkin's disease, childhood
C0279921|T191|NSHD, childhood
C0279921|T191|NS HD, childhood
C0279921|T191|HD, nodular sclerosis, childhood
C0279921|T191|lymphoma, nodular sclerosing childhood Hodgkin's
C1334425|T191|Low Grade Malignant Neoplasm
C0449443|T034|Receptor Status
C0449443|T034|Receptor status
C0449443|T034|Receptor status (attribute)
C0862640|T191|Stage I Prostate Adenocarcinoma
C0862640|T191|Stage I Prostate Adenocarcinoma AJCC v7
C116432|T061|Image-Guided Adaptive Radiation Therapy
C0278861|T191|Recurrent Thyroid Gland Carcinoma
C0278861|T191|Recurrent Cancer of Thyroid Gland
C0278861|T191|Recurrent Thyroid Carcinoma
C0278861|T191|Recurrent Cancer of Thyroid
C0278861|T191|thyroid cancer, recurrent
C0278861|T191|Relapsed Cancer of the Thyroid Gland
C0278861|T191|Relapsed Cancer of Thyroid Gland
C0278861|T191|Relapsed Cancer of the Thyroid
C0278861|T191|Recurrent Cancer of the Thyroid Gland
C0278861|T191|Recurrent Cancer of the Thyroid
C0278861|T191|Relapsed Thyroid Gland Cancer
C0278861|T191|recurrent thyroid cancer
C0278861|T191|Thyroid cancer recurrent
C0278861|T191|Recurrent Thyroid Cancer
C0278861|T191|Relapsed Thyroid Cancer
C0278861|T191|Relapsed Cancer of Thyroid
C1333851|T191|Grade 3b Malignant Neoplasm
C0085533|T061|Adjuvant Chemotherapy
C0085533|T061|DRUG THER ADJUVANT
C0085533|T061|CHEMOTHER ADJUVANT
C0085533|T061|ADJUVANT DRUG THER
C0085533|T061|Chemotherapy, Adjuvant
C0085533|T061|Drug Therapy, Adjuvant
C0085533|T061|Adjuvant Drug Therapy
C1275387|T201|Tumor size after sectioning
C1275387|T201|Tumour dimension after sectioning
C1275387|T201|Tumor size after sectioning (observable entity)
C1275387|T201|Tumour size after sectioning
C1275387|T201|Tumor dimension after sectioning
C1709447|T191|Paget Disease of the Breast without Invasive Carcinoma
C1709447|T191|Paget's Disease of the Breast without Invasive Carcinoma
C1709447|T191|Tis (Paget)
C1321210|T033|Tumor nodule size, greatest dimension
C1321210|T033|Tumor nodule size, greatest dimension (observable entity)
C1321210|T033|Tumour nodule size, greatest dimension
C0280402|T191|Recurrent Laryngeal Verrucous Carcinoma
C0280402|T191|Recurrent Verrucous Carcinoma of the Larynx
C0280402|T191|Relapsed Verrucous Carcinoma of the Larynx
C0280402|T191|Relapsed Laryngeal Verrucous Carcinoma
C0280402|T191|Relapsed Larynx Verrucous Carcinoma
C0280402|T191|Laryngeal verrucous carcinoma recurrent
C0280402|T191|recurrent verrucous carcinoma of the larynx
C0280402|T191|larynx verrucous carcinoma, recurrent
C0280402|T191|Relapsed Verrucous Carcinoma of Larynx
C0280402|T191|Recurrent Larynx Verrucous Carcinoma
C0280402|T191|verrucous carcinoma of the larynx, recurrent
C0280402|T191|laryngeal verrucous carcinoma, recurrent
C0280402|T191|Recurrent Verrucous Carcinoma of Larynx
C1333845|T191|Grade 3 Malignant Neoplasm
C0281464|T191|AIDS-Related Lymphoblastic Lymphoma
C0281464|T191|AIDS Related Lymphoblastic lymphoma
C0281464|T191|AIDS Associated Lymphoblastic lymphoma
C0281464|T191|AIDS-Associated Lymphoblastic lymphoma
C0281464|T191|AIDS-Related Precursor Lymphoblastic Lymphoma
C1515863|T191|Acinar Prostate Adenocarcinoma, Foamy Gland Variant
C0742078|T047|Brain Mass
C0742078|T047|Space-occupying lesion of brain
C0742078|T047|Mass lesion of brain (finding)
C0742078|T047|Brain mass
C0742078|T047|Mass lesion of brain
C0085203|T061|Stereotactic Radiosurgery
C0085203|T061|stereotaxic radiation therapy
C0085203|T061|STEREOTACTIC RADIOSURG
C0085203|T061|Stereo radiosurgery NOS
C0085203|T061|Stereotactic radiosurgery (procedure)
C0085203|T061|Stereotactic Radiotherapy
C0085203|T061|SBRT
C0085203|T061|Radiosurgeries
C0085203|T061|Radiosurgery
C0085203|T061|Stereotactic External Beam Irradiation
C0085203|T061|Radiosurgery, Stereotactic
C0085203|T061|RADIOSURG STEREOTACTIC
C0085203|T061|stereotaxic radiosurgery
C0085203|T061|Stereotactic Radiation Therapy
C0085203|T061|Stereotactic radiosurgery, not otherwise specified
C0085203|T061|stereotactic body radiation therapy
C0085203|T061|RADIOSURG
C0085203|T061|Stereotactic radiosurgery
C0085203|T061|Radiosurgeries, Stereotactic
C0085203|T061|Stereotactic Radiosurgeries
C0085203|T061|stereotactic radiation therapy
C0085203|T061|stereotactic radiosurgery
C0085203|T061|stereotactic external-beam radiation therapy
C0854762|T191|Recurrent Esophageal Adenocarcinoma
C0854762|T191|Oesophageal adenocarcinoma recurrent
C0854762|T191|Recurrent Adenocarcinoma of the Esophagus
C0854762|T191|Relapsed Adenocarcinoma of the Esophagus
C0854762|T191|Esophageal adenocarcinoma recurrent
C0854762|T191|Oesophageal Adenocarcinoma Recurrent
C0854762|T191|Esophageal Adenocarcinoma, Recurrent
C0854762|T191|Relapsed Esophagus Adenocarcinoma
C0854762|T191|Recurrent Esophagus Adenocarcinoma
C0854762|T191|Relapsed Adenocarcinoma of Esophagus
C0854762|T191|Recurrent Adenocarcinoma of Esophagus
C0854762|T191|Relapsed Esophageal Adenocarcinoma
C0746765|T033|Nasal Mass
C0746765|T033|Mass of Nose
C0746765|T033|Mass of nose (finding)
C0746765|T033|Mass of nose
C0746765|T033|Mass of the Nose
CL433924|T191|Recurrent Childhood Anaplastic Oligodendroglioma
CL433924|T191|recurrent childhood anaplastic oligodendroglioma
C0238736|T033|Mass of the Back
C0238736|T033|Mass of Back
C0279920|T191|Childhood Lymphocyte Depleted Classical Hodgkin Lymphoma
C0279920|T191|Childhood Lymphocyte Depleted Hodgkin Lymphoma
C0279920|T191|childhood lymphocyte depletion Hodgkin lymphoma
C0279920|T191|childhood HD, lymphocyte depletion
C0279920|T191|Childhood Lymphocyte Depleted Hodgkin's Lymphoma
C0279920|T191|Pediatric Lymphocyte Depleted Hodgkin's Lymphoma
C0279920|T191|HDLD, childhood
C0279920|T191|pediatric HD, lymphocyte depletion
C0279920|T191|pediatric Hodgkin's disease, lymphocyte depletion
C0279920|T191|lymphoma, lymphocyte depleted childhood Hodgkin's
C0279920|T191|childhood lymphocyte depletion Hodgkin's disease
C0279920|T191|Childhood LDHD
C0279920|T191|LDHD, childhood
C0279920|T191|childhood Hodgkin's disease, lymphocyte depleted
C0279920|T191|Hodgkin's disease, lymphocyte depleted, childhood
C0279920|T191|Childhood Lymphocyte Depletion Hodgkin's Disease
C0279920|T191|lymphocyte depleted Hodgkin's disease, childhood
C0279920|T191|LD HD, childhood
C0279920|T191|Pediatric Lymphocyte Depletion Hodgkin's Lymphoma
C0279920|T191|pediatric lymphocyte depletion Hodgkin's disease
C0279920|T191|Pediatric LDHD
C0279920|T191|HD LD, childhood
C0279920|T191|lymphocyte depleted HD, childhood
C0279920|T191|lymphocyte depletion Hodgkin's disease, childhood
C0279920|T191|Childhood Lymphocyte Depletion Hodgkin's Lymphoma
C0279920|T191|lymphocyte depletion HD, childhood
C0279920|T191|HD lymphocyte depleted, childhood
C0279920|T191|Pediatric Lymphocyte Depletion Hodgkin's Disease
C1335717|T191|Recurrent Non-Cutaneous Melanoma
C1332216|T191|Adult Systemic Anaplastic Large Cell Lymphoma
C1332216|T191|Adult Systemic CD30+ Anaplastic Large Cell Lymphoma
C1332216|T191|Adult Systemic K-1+ Anaplastic Large Cell Lymphoma
C0544885|T049|Nonsense Mutation
C0544885|T049|Nonsense mutation (finding)
C0544885|T049|Premature Termination Abnormality
C0544885|T049|nonsense mutation
C0544885|T049|Nonsense Mutations
C0544885|T049|Premature Termination Mutation
C0544885|T049|Nonsense mutation
C0544885|T049|Mutation, Nonsense
C0544885|T049|Mutations, Nonsense
C0024886|T061|Total Mastectomy
C0024886|T061|Mastectomies, Total
C0024886|T061|Unilateral Mastectomy, complete
C0024886|T061|Unilateral mastectomy (situation)
C0024886|T061|Unilateral simple mastectomy (situation)
C0024886|T061|SM - Simple mastectomy
C0024886|T061|Simple mastectomy (procedure)
C0024886|T061|Mastectomies, Simple
C0024886|T061|Total mastectomy
C0024886|T061|Simple Mastectomy
C0024886|T061|Unilat simple mastectomy
C0024886|T061|Unilateral simple mastectomy
C0024886|T061|simple mastectomy
C0024886|T061|total mastectomy
C0024886|T061|Simple Mastectomies
C0024886|T061|Unilateral Mastectomy, NOS
C0024886|T061|Total Mastectomies
C0024886|T061|Mastectomy, Simple
C0024886|T061|Mastectomy, Total
C0024886|T061|Unilateral mastectomy
C0024886|T061|Simple mastectomy
C0024886|T061|Mastectomy
C1883168|T061|Stationary Beam Radiation Therapy
C1883168|T061|Fixed Beam Radiation Therapy
C1883168|T061|Fixed Beam
C1883168|T061|Stationary Beam Radiation
C1883168|T061|Fixed Beam Radiation
C1336814|T191|Transplant-Related Malignant Neoplasm
C1336814|T191|Transplant-Related Cancer
C1336814|T191|Transplant-Related Malignancy
C0280182|T191|Recurrent Grade 1 Follicular Lymphoma
C0280182|T191|follicular small cleaved cell lymphoma, recurrent
C0280182|T191|Relapsed Grade I Follicular Small Cleaved Cell Lymphoma
C0280182|T191|recurrent grade I follicular small cleaved cell lymphoma
C0280182|T191|Recurrent Grade I Follicular Small Cleaved Cell Lymphoma
C0280182|T191|Recurrent Follicular Small Cleaved Cell Lymphoma
C0280182|T191|Recurrent Grade I Follicular Lymphoma
C0280182|T191|follicular small cleaved cell lymphoma, relapsed
C0280182|T191|recurrent grade 1 follicular lymphoma
C0280182|T191|relapsed follicular small cleaved cell lymphoma
C0280182|T191|Relapsed Follicular Small Cleaved Cell Lymphoma
C0280182|T191|Relapsed Grade I Follicular Lymphoma
C0854747|T191|Stage IV AIDS-Related Anal Canal Cancer
C0854747|T191|Stage IV AIDS-Related Anal Canal Cancer AJCC v7
C0854747|T191|Stage IV AIDS-Related Anal Canal Cancer AJCC v6
C1710404|T049|Thymidine to Adenosine Transversion Abnormality
C1710404|T049|Thymidine to Adenosine Mutation
C1710404|T049|Thymidine to Adenosine Transversion
C0935916|T121|Fulvestrant
C0935916|T121|ZD9238
C0935916|T121|ICI 182780
C0935916|T121|7a-[9-[(4,4,5,5,5,-Pentafluoropentyl)sulphinyl]nonyl]-estra-1,3,5(10)-triene-3,17b-diol
C0935916|T121|Faslodex(ICI 182,780)
C0935916|T121|FULVESTRANT
C0935916|T121|Faslodex
C0935916|T121|fulvestrant
C0935916|T121|ICI 182,780
CL446011|T061|Scattering Proton Beam Therapy
C0280366|T191|Recurrent Oral Cavity Mucoepidermoid Carcinoma
C0280366|T191|Relapsed Oral Cavity Mucoepidermoid Carcinoma
C0280366|T191|Mucoepidermoid carcinoma of the oral cavity recurrent
C0280366|T191|Recurrent Mucoepidermoid Carcinoma of the Oral Cavity
C0280366|T191|Recurrent Mouth Mucoepidermoid Carcinoma
C0280366|T191|Recurrent Mucoepidermoid Carcinoma of Oral Cavity
C0280366|T191|Relapsed Mucoepidermoid Carcinoma of the Oral Cavity
C0280366|T191|Relapsed Mucoepidermoid Carcinoma of Mouth
C0280366|T191|Relapsed Mucoepidermoid Carcinoma of the Mouth
C0280366|T191|oral cavity mucoepidermoid carcinoma, recurrent
C0280366|T191|Relapsed Mucoepidermoid Carcinoma of Oral Cavity
C0280366|T191|recurrent mucoepidermoid carcinoma of the oral cavity
C0280366|T191|mucoepidermoid carcinoma of the oral cavity, recurrent
C0280366|T191|Relapsed Mouth Mucoepidermoid Carcinoma
C0280366|T191|Recurrent Mucoepidermoid Carcinoma of the Mouth
C0280366|T191|Recurrent Mucoepidermoid Carcinoma of Mouth
C0278735|T191|Stage I Childhood Lymphoblastic Lymphoma
C0278735|T191|Pediatric Lymphoblastic Lymphoma Stage I
C0278735|T191|Stage I Childhood Precursor Lymphoblastic Lymphoma
C0278735|T191|Childhood Lymphoblastic Lymphoma Stage I
C0278735|T191|Stage I Pediatric Lymphoblastic Lymphoma
C2825183|T061|Ventricular Ablation
C2825183|T061|ABLATION, VENTRICULAR
C056507|T114|Gemcitabine
C056507|T114|2,2 difluorodexoycytidine
C056507|T114|gemcitabine [Chemical/Ingredient]
C056507|T114|1-(2-Oxo-4-amino-1,2-dihydropyrimidin-1-yl)-2-deoxy-2,2-difluororibose
C056507|T114|gemcitabine
C056507|T114|613327
C056507|T114|2'-deoxy-2'-difluorocytidine
C056507|T114|2',2'-difluorodeoxycytidine
C056507|T114|47762
C056507|T114|Gemcitabine (substance)
C056507|T114|GEMCITABINE
C056507|T114|2',2'-DFDC
C056507|T114|2',2'-difluoro-2'-deoxycytidine
C056507|T114|103882-84-4
C056507|T114|Gemcitabine (product)
C056507|T114|Difluorodeoxycytidine
C056507|T114|dFdC
C056507|T114|2'Deoxy-2',2'-Difluorocytidine
C056507|T114|dFdCyd
C2986679|T191|Stage III Childhood Non-Hodgkin Lymphoma
C2986679|T191|stage III childhood non-Hodgkin lymphoma
C1334574|T191|Malignant Childhood Germ Cell Tumor
C1334574|T191|Malignant Pediatric Germ Cell Neoplasm
C1334574|T191|Malignant Childhood Germ Cell Neoplasm
C1334574|T191|Malignant Pediatric Germ Cell Tumor
C0239059|T131|Cigarette Smoking
C0239059|T131|Cigarette smoke (substance)
C0239059|T131|Cigarette smoking behavior
C0239059|T131|CIGARETTE SMOKING
C0239059|T131|Cigarette smoking
C0239059|T131|Smoking, Cigarette
C0239059|T131|cigarette smoking
C0239059|T131|Cigarette smoke
C0204032|T061|Infrared Radiation Therapy
C0204032|T061|infrared radiation therapy
C0204032|T061|Radiant heat: infrared:physio.
C0204032|T061|Infrared therapy
C0204032|T061|Radiant heat therapy
C0204032|T061|Infrared radiation therapy (regime/therapy)
C0204032|T061|Infrared radiation therapy
C1332222|T191|Aflatoxins-Related Hepatocellular Carcinoma
C0013089|T121|Doxorubicin
C0013089|T121|Doxorubicin (substance)
C0013089|T121|14-hydroxydaunorubicine
C0013089|T121|Hydroxyl Daunorubicin
C0013089|T121|5,12-Naphthacenedione, 10-((3-amino-2,3,6-trideoxy-alpha-L-lyxo-hexopyranosyl)oxy)-7,8,9,10-tetrahydro-6,8,11-trihydroxy-8-(hydroxyacetyl)-1-methoxy-, (8S-cis)-
C0013089|T121|Doxorubicin [Chemical/Ingredient]
C0013089|T121|adriamycin
C0013089|T121|14-Hydroxydaunomycin
C0013089|T121|Hydroxyldaunorubicin
C0013089|T121|DOXOrubicin
C0013089|T121|DOXORUBICIN
C0013089|T121|doxorubicin
C0013089|T121|(8S-cis)-10-[(3-Amino-2,3,6-trideoxy-alpha-L-lyxo-hexopyranosyl)oxy]-7,8,9,10-tetrahydro-6,8,11-trihydroxy-8-(hydroxyacetyl)-1-methoxy-5,12-naphthacenedione
C0013089|T121|(8S-cis)-10-[(3-Amino-2,3,6-trideoxy-alpha-L-lyxo-hexopyranosyl)oxy]-7,8,9,10-tetrahydro-6,8,11-trihydroxy-8-(hydroacetyl)-1-methoxy-5,12-naphthacenedione
C0013089|T121|Doxorubicin (product)
C2986611|T033|Dirty Necrosis
C2986611|T033|dirty necrosis
C1332078|T191|Anaplastic Large Cell Lymphoma, ALK-Negative
C1332078|T191|ALK-Negative Anaplastic Large Cell Lymphoma
C1332078|T191|ALCL, ALK-
C0085101|T061|Radioimmunotherapy
C0085101|T061|radioimmunotherapy
C0085101|T061|RADIOIMMUNOTHER
C0085101|T061|Immunoradiotherapy
C0085101|T061|radioimmunotherapeutics
C0085101|T061|Immunoradiotherapies
C0085101|T061|Radioimmunotherapy (procedure)
C0085101|T061|Radioimmunotherapies
C0085101|T061|IMMUNORADIOTHER
C0085101|T061|Immunotherapy, Cancer, Radioisotope
C114968|T191|Childhood Gliosarcoma
C114968|T191|childhood gliosarcoma
C1332643|T191|Burkitt Lymphoma Post-Transplant Lymphoproliferative Disorder
C1332643|T191|Burkitt's Lymphoma Post-Transplant Lymphoproliferative Disorder
C1332643|T191|Burkitt Lymphoma PTLD
C1332643|T191|Burkitt's Lymphoma PTLD
C0853972|T191|Stage IV Inflammatory Breast Carcinoma
C0853972|T191|Stage IV Inflammatory Breast Cancer
C0853972|T191|Inflammatory Carcinoma of Breast Stage IV
C0278716|T191|Recurrent Renal Wilms Tumor
C0278716|T191|Recurrent Kidney Adenosarcoma
C0278716|T191|nephroblastoma, recurrent
C0278716|T191|recurrent Wilms tumor
C0278716|T191|Recurrent Renal Adenosarcoma
C0278716|T191|recurrent Wilm's tumor
C0278716|T191|Wilm's tumor, recurrent
C0278716|T191|Recurrent Nephroblastoma
C0278716|T191|recurrent nephroblastoma
C0278716|T191|Relapsed Renal Adenosarcoma
C0278716|T191|Relapsed Nephroblastoma
C0278716|T191|Wilms tumor, recurrent
C0278716|T191|Relapsed Kidney Adenosarcoma
C0278716|T191|Wilms' tumor, recurrent
C0278716|T191|Recurrent Renal Wilms' Tumor
C0278716|T191|Relapsed Renal Wilms' Tumor
C1333126|T033|Comedo Necrosis
C1333126|T033|Comedo Change
C1333126|T033|Comedo Lesion
C1333126|T033|Comedo-Like Necrosis
C0861727|T191|Metastatic Pancreatic Adenocarcinoma
C0861727|T191|Pancreatic adenocarcinoma metastatic
C0677725|T191|Recurrent Mantle Cell Lymphoma
C0677725|T191|recurrent mantle cell lymphoma
C0677725|T191|Mantle cell lymphoma recurrent
C0278812|T191|Recurrent Extrahepatic Bile Duct Carcinoma
C0278812|T191|Recurrent Extrahepatic Bile Duct Cancer
C0278812|T191|Recurrent Cancer of Extrahepatic Bile Duct
C0278812|T191|Relapsed Cancer of Extrahepatic Bile Duct
C0278812|T191|Relapsed Cancer of the Extrahepatic Bile Duct
C0278812|T191|bile duct cancer, recurrent extrahepatic
C0278812|T191|extrahepatic bile duct cancer, recurrent
C0278812|T191|recurrent extrahepatic bile duct cancer
C0278812|T191|Recurrent Cancer of the Extrahepatic Bile Duct
CL448216|T191|Metastatic Malignant Neoplasm to the Ovary
CL448216|T191|Metastatic Malignant Tumor to the Ovary
CL448216|T191|Metastases to Ovary
CL448216|T191|Ovarian Metastasis
CL448216|T191|Metastasis to Ovary
C2986508|T061|Unsealed Internal Radiation Therapy
C2986508|T061|unsealed internal radiation therapy
C1300494|T201|Tumor size, dominant nodule, greatest dimension
C1300494|T201|Tumour size, dominant nodule, greatest dimension
C1300494|T201|Tumor size, dominant nodule, greatest dimension (observable entity)
C3273217|T191|Invasive Lobular Breast Carcinoma, Solid Variant
C0220621|T191|Childhood Acute Myeloid Leukemia
C0220621|T191|acute myeloid leukemia, childhood
C0220621|T191|Childhood Acute Myelocytic Leukemia
C0220621|T191|childhood acute myelogenous leukemia
C0220621|T191|acute myeloblastic leukemia, childhood
C0220621|T191|childhood leukemia, acute myelogenous
C0220621|T191|Pediatric AML
C0220621|T191|AML, childhood
C0220621|T191|pediatric leukemia, acute myeloid
C0220621|T191|childhood acute granulocytic leukemia
C0220621|T191|leukemia, pediatric acute myelogenous
C0220621|T191|pediatric acute granulocytic leukemia
C0220621|T191|AGL, pediatric
C0220621|T191|leukemia, childhood acute myelogenous
C0220621|T191|AML, pediatric
C0220621|T191|Pediatric Acute Myelocytic Leukemia
C0220621|T191|leukemia, pediatric acute myeloid
C0220621|T191|childhood acute myelocytic leukemia
C0220621|T191|myeloid leukemia, pediatric acute
C0220621|T191|acute myelogenous leukemia, childhood
C0220621|T191|acute myelocytic leukemia, childhood
C0220621|T191|acute myeloid leukemia, pediatric
C0220621|T191|acute myelogenous leukemia, pediatric
C0220621|T191|granulocytic leukemia, childhood acute
C0220621|T191|leukemia, childhood acute myeloblastic
C0220621|T191|AGL, childhood
C0220621|T191|pediatric AGL
C0220621|T191|Childhood AML
C0220621|T191|pediatric leukemia, acute myelogenous
C0220621|T191|acute granulocytic leukemia, childhood
C0220621|T191|Acute myeloid leukemia (AML), child
C0220621|T191|Childhood Acute Myeloblastic Leukemia
C0220621|T191|Childhood Acute Granulocytic Leukemia
C0220621|T191|pediatric acute myeloid leukemia
C0220621|T191|Pediatric Acute Myelogenous Leukemia
C0220621|T191|myelogenous leukemia, pediatric acute
C0220621|T191|Pediatric Acute Myeloblastic Leukemia
C0220621|T191|childhood AML
C0220621|T191|pediatric acute myelogenous leukemia
C0220621|T191|myeloblastic leukemia, childhood acute
C0220621|T191|leukemia, childhood acute myeloid
C0220621|T191|childhood acute myeloblastic leukemia
C0220621|T191|pediatric acute myeloblastic leukemia
C0220621|T191|Pediatric Acute Myeloid Leukemia
C0220621|T191|Leukemia, acute myeloid (AML), child
C0220621|T191|myelocytic leukemia, childhood acute
C0220621|T191|pediatric acute myelocytic leukemia
C0220621|T191|pediatric AML
C0220621|T191|myeloid leukemia, childhood acute
C0220621|T191|childhood leukemia, acute myeloid
C0220621|T191|myelogenous leukemia, childhood acute
C0220621|T191|Childhood Acute Myelogenous Leukemia
C0333513|T046|Fibrinoid Necrosis
C0333513|T046|fibrinoid degeneration (morphologic abnormality)
C0333513|T046|fibrinoid degeneration
C0333513|T046|Fibrinoid necrosis
C0333513|T046|Fibrinoid necrosis (morphologic abnormality)
C0333513|T046|Fibrinoid degeneration
C0280790|T191|Adult Anaplastic Oligodendroglioma
C0280790|T191|anaplastic oligodendroglioma, adult
C0280790|T191|Adult Undifferentiated Oligodendroglioma
C0280790|T191|oligodendroglioma, adult anaplastic
C0280790|T191|adult anaplastic oligodendroglioma
C0879257|T191|Hereditary Papillary Renal Cell Carcinoma
C0879257|T191|Hereditary Papillary Carcinoma of Kidney
C0879257|T191|Hereditary Papillary Renal Carcinoma
C0879257|T191|hereditary papillary renal cell carcinoma
C0879257|T191|Hereditary papillary renal carcinoma
C0879257|T191|Hereditary Papillary Carcinoma of the Kidney
C0879257|T191|Hereditary Kidney Papillary Carcinoma
C0879257|T191|Familial Renal Papillary Carcinoma
CL414683|T191|Metastatic Carcinoma to the Bone
CL414683|T191|Bone Carcinoma
C1301451|T201|Maximum thickness of diffuse tumor
C1301451|T201|Maximum thickness of diffuse tumour
C1301451|T201|Maximum thickness of diffuse tumor (observable entity)
C1516076|T033|Asymptomatic Mass
C0497565|T191|Malignant Neoplasm
C0497565|T191|Neoplasm, malignant
C0497565|T191|Malignant Nervous System Neoplasm
C0497565|T191|MALIGNANCY
C0497565|T191|Cancer (NOS)
C0497565|T191|Unclassified tumour, malignant
C0497565|T191|Tumor, malignant
C0497565|T191|CANCER (NOS)
C0497565|T191|Cancers
C0497565|T191|Malignant Nervous System Tumor
C0497565|T191|Tumour, malignant
C0497565|T191|malignant neoplastic disease
C0497565|T191|Malignant neoplasms (C00-C96)
C0497565|T191|Cancer NOS
C0497565|T191|malignant neurologic neoplasms
C0497565|T191|Neoplasm malignant
C0497565|T191|cancer
C0497565|T191|Malignant obstetric neoplasm
C0497565|T191|Malignant neoplastic disease
C0497565|T191|Primary Malignant Neoplasm
C0497565|T191|Malignant neoplasm of nervous system
C0497565|T191|Malignant Neoplastic Disease
C0497565|T191|Malignant tumour of nervous system
C0497565|T191|Malignant tumour morphology
C0497565|T191|Malignant neoplasm, primary (morphologic abnormality)
C0497565|T191|Blastoma
C0497565|T191|Malignant tumor morphology
C0497565|T191|Cancer
C0497565|T191|CA - Cancer
C0497565|T191|Malignant Neoplasms
C0497565|T191|Malignant tumour
C0497565|T191|Malignant Neoplasm of Nervous System
C0497565|T191|NEOPLASM, MALIGNANT
C0497565|T191|malignant neoplasm
C0497565|T191|Neoplasm, malignant (primary)
C0497565|T191|Malignancy
C0497565|T191|Cancer morphology
C0497565|T191|Malignant neoplasm NOS
C0497565|T191|Malignant neoplasm of nervous system NOS
C0497565|T191|Malignant tumor
C0497565|T191|Malignant neoplasm, unspecified
C0497565|T191|Malignancy, unspecified site
C0497565|T191|neoplasm/cancer
C0497565|T191|Primary malignant neoplasm
C0497565|T191|Malignant neoplasm
C0497565|T191|MALIGNANT NEOPLASM
C0497565|T191|malignant tumor
C0497565|T191|Primary malignant neoplasm (disorder)
C0497565|T191|CANCER
C0497565|T191|Nervous System Neoplasms, Malignant
C0497565|T191|Malignant Tumor
C0497565|T191|NEOPLASM MALIGNANT
C0497565|T191|Malignant neoplasm of nervous system (disorder)
C0497565|T191|Malignant neurologic neoplasms
C0497565|T191|Malignant nervous system neoplasm
C0497565|T191|CA
C0497565|T191|Cancer, unspecified site
C0497565|T191|MALIGNANT TUMOR
C0497565|T191|Malignant neoplasm without specification of site
C0497565|T191|Malignant neoplastic disease (disorder)
C0497565|T191|Malignant neoplasms
C0497565|T191|Malignant nervous system neoplasm NOS
C0497565|T191|Malignant tumor of nervous system
C0497565|T191|Malignant Tumor of Nervous System
C0497565|T191|Malignant Tumor of the Nervous System
C0497565|T191|MALIGNANCIES
C0497565|T191|Malignant Neoplasm of the Nervous System
C0497565|T191|Malignant neoplasm, primary
C0497565|T191|malignancy
C0497565|T191|Unclassified tumor, malignant
C0497565|T191|malignant tumoral disease
C0497565|T191|Tumor, malignant, NOS
C0279085|T191|Kaposi Sarcoma Related to Immunosuppressive Treatment
C0279085|T191|Kaposi's Sarcoma Related to Immunosuppressive Treatment
C0279085|T191|Immunosuppressive Treatment Related Kaposi Sarcoma
C0279085|T191|Immunosuppressive Treatment Related Kaposi's Sarcoma
C0279564|T191|Invasive Lobular Breast Carcinoma with Predominant In Situ Component
C0279564|T191|Infiltrating Lobular Breast Carcinoma with Predominant In Situ Component
C0085090|T191|AIDS-Related Lymphoma
C0085090|T191|AIDS Lymphoma
C0085090|T191|Lymphoma AIDS Related
C0085090|T191|HIV Associated Lymphoma
C0085090|T191|Lymphoma, AIDS-Related
C0085090|T191|AIDS Related Lymphoma
C1332235|T191|Alkylating Agent-Related Myelodysplastic Syndrome
C1332235|T191|Alkylating Agent Related Myelodysplastic Syndrome
C1334157|T191|Immunoblastic Lymphoma Post-Transplant Lymphoproliferative Disorder
C1334157|T191|Immunoblastic Lymphoma PTLD
C1334157|T191|Immunoblastic Diffuse Large B-Cell Lymphoma PTLD
CL415252|T191|Recurrent Hepatocellular Carcinoma
CL415252|T191|Relapsed Carcinoma of the Liver Cell
CL415252|T191|Hepatocellular carcinoma recurrent
CL415252|T191|Relapsed Carcinoma of Liver Cell
CL415252|T191|Hepatocellular Carcinoma, Recurrent
CL415252|T191|Recurrent Liver Cell Carcinoma
CL415252|T191|Recurrent Hepatoma
CL415252|T191|Recurrent Carcinoma of Liver Cell
CL415252|T191|Relapsed Hepatocellular Carcinoma
CL415252|T191|Hepatoma recurrent
CL415252|T191|Relapsed Liver Cell Carcinoma
CL415252|T191|Relapsed Hepatoma
CL415252|T191|Recurrent Carcinoma of the Liver Cell
CL472494|T191|Childhood Central Nervous System Embryonal Neoplasm
C1334749|T191|Methotrexate-Associated Lymphoproliferative Disorder
C1334749|T191|Methotrexate-Associated Lymphoproliferation
C1332978|T191|Childhood Lymphocyte-Rich Classical Hodgkin Lymphoma
C1332978|T191|Childhood Lymphocyte Rich Classical Hodgkin's Lymphoma
C1332978|T191|Childhood Lymphocyte Rich Classical Hodgkin's Disease
C1332978|T191|Pediatric Lymphocyte Rich Classical Hodgkin's Lymphoma
C1332978|T191|Childhood Lymphocyte Rich Classical Hodgkin Lymphoma
C1332978|T191|Pediatric Lymphocyte Rich Classical Hodgkin's Disease
C0281241|T191|AIDS-Related Primary Central Nervous System Lymphoma
C0281241|T191|AIDS-Related Primary CNS Lymphoma
C0281241|T191|AIDS-Related Lymphoma of Primary Central Nervous System
C0281241|T191|AIDS Related Primary Central Nervous System Lymphoma
C0281241|T191|AIDS Related Lymphoma of the Primary Central Nervous System
C0281241|T191|AIDS Related Lymphoma of Primary Central Nervous System
C0281241|T191|AIDS-related primary CNS lymphoma
C0281241|T191|AIDS-Related Lymphoma of the Primary Central Nervous System
C0281241|T191|AIDS Related Primary CNS Lymphoma
C114451|T191|Rare Malignant Childhood Neoplasm
C115030|T191|Stage II Childhood Anaplastic Large Cell Lymphoma
C0346973|T191|Metastatic Malignant Neoplasm to the Large Intestine
C0346973|T191|Metastases to Large Intestine
C0346973|T191|Metastatic Tumor to the Large Intestine
C0346973|T191|Metastasis to the Large Bowel
C0346973|T191|Metastasis to Large Bowel
C0346973|T191|Metastatic Neoplasm to the Large Intestine
C0346973|T191|Metastasis to the Large Intestine
C1512739|T191|Infiltrating Bladder Urothelial Carcinoma, Lymphoma-Like Variant
C0014582|T121|Epirubicin
C0014582|T121|IMI 28
C0014582|T121|4'-Epiadriamycin
C0014582|T121|Epirubicin (product)
C0014582|T121|EPIRUBICIN
C0014582|T121|epi DX
C0014582|T121|EPIADRIAMYCIN 04
C0014582|T121|4'-Epidoxorubicin
C0014582|T121|(8S-cis)-10-((3-Amino-2,3,6-trideoxy-beta-L-arabino-hexopyranosyl)oxy)-7,8,9,10-tetrahydro-6,8,11-trihydroxy-8-(hydroxyacetyl)-1-methoxy-5,12-naphthacenedione
C0014582|T121|pidorubicin
C0014582|T121|epidoxorubicin
C0014582|T121|4' Epidoxorubicin
C0014582|T121|Epi DX
C0014582|T121|4'-epi-doxorubicin
C0014582|T121|Epirubicin [Chemical/Ingredient]
C0014582|T121|4'-epi-adriamycin
C0014582|T121|3-Glycoloyl-1,2,3,4,6,11-hexahydro-3,5,12-trihydroxy-10-methoxy-6,11-dioxo-1-naphthacenyl-3-amino-2,3,6-trideoxy-alpha-L-arabino-hexopyranoside
C0014582|T121|4' Epiadriamycin
C0014582|T121|Pidorubicin
C0014582|T121|4' Epi Adriamycin
C0014582|T121|4' Epi DXR
C0014582|T121|4'-epidoxorubicin
C0014582|T121|4'-epi-DX
C0014582|T121|4'-Epi-Doxorubicin
C0014582|T121|4'-Epi-DXR
C0014582|T121|4' Epi Doxorubicin
C0014582|T121|4'-epi DX
C0014582|T121|IMI28
C0014582|T121|4'-Epi-Adriamycin
C0014582|T121|Epidoxorubicin
C0014582|T121|EPIDOXORUBICIN 04
C0014582|T121|5,12-Naphthacenedione, 10-((3-amino-2,3,6-trideoxy-alpha-L-arabino-hexopyranosyl)oxy)-7,8,9,10-tetrahydro-6,8,11-trihydroxy-8-(hydroxyacetyl)-1-methoxy-, (8S-cis)-
C0014582|T121|epirubicin
C0014582|T121|Epirubicin (substance)
C0014582|T121|IMI-28
C0014582|T121|epi-ADR
C0014582|T121|4'-epiadriamycin
C0686112|T191|Metastatic Malignant Neoplasm to the Gallbladder
C0686112|T191|Metastatic Tumor to the Gallbladder
C0686112|T191|Secondary Malignant Neoplasm to the Gallbladder
C0686112|T191|Metastatic Neoplasm to the Gallbladder
C0686112|T191|Secondary Malignant Tumor to the Gallbladder
C0206624|T191|Hepatoblastoma
C0206624|T191|Malignant neoplasm: Hepatoblastoma
C0206624|T191|childhood hepatoblastoma
C0206624|T191|Hepatoblastoma (disorder)
C0206624|T191|pediatric hepatoblastoma
C0206624|T191|Pediatric Embryonal Hepatoma
C0206624|T191|Hepatoblastoma (clinical)
C0206624|T191|PEDIATRIC HEPATOBLASTOMA
C0206624|T191|HBL - Hepatoblastoma
C0206624|T191|HBL
C0206624|T191|Pediatric Hepatoblastoma
C0206624|T191|Hepatoblastoma (morphologic abnormality)
C0206624|T191|hepatoblastoma, childhood
C0206624|T191|Embryonal hepatoma
C0206624|T191|PEDIATRIC EMBRYONAL HEPATOMA
C0206624|T191|Hepatoblastomas
C0206624|T191|Hepatoblastoma NOS
C0206624|T191|HEPATOBLASTOMA
C0206624|T191|hepatoblastoma
C0206624|T191|Hepatoblastoma [Disease/Finding]
C0206624|T191|HEPATOBLASTOMA, MALIGNANT
C0206624|T191|Hepatoblastoma of liver
C0280745|T191|Secondary Myelodysplastic Syndrome
C0280745|T191|secondary myelodysplastic syndrome
C0280745|T191|Secondary MDS
C0280745|T191|secondary myelodysplastic syndromes
C0280745|T191|secondary MDS
C0280745|T191|myelodysplastic syndromes, secondary
C1709092|T049|Multiple Nucleotide Abnormalities
CL448282|T191|Recurrent Nasal Type NK/T-Cell Lymphoma
CL448282|T191|Recurrent Angiocentric Lymphoma
CL448282|T191|Relapsed Angiocentric Lymphoma
CL448282|T191|Relapsed Nasal Type NK/T-Cell Lymphoma
C1512742|T191|Infiltrating Bladder Urothelial Carcinoma, Plasmacytoid Variant
C0279016|T061|Low-LET Electron Therapy
C1332953|T191|Childhood Central Nervous System Germinoma
C1332953|T191|childhood central nervous system germinoma
C1332953|T191|childhood CNS germinoma
C0278818|T191|Recurrent Adrenal Cortex Carcinoma
C0278818|T191|Recurrent Carcinoma of the Adrenal Cortex
C0278818|T191|Relapsed Adrenocortical Carcinoma
C0278818|T191|adrenocortical carcinoma, recurrent
C0278818|T191|Relapsed Carcinoma of the Adrenal Cortex
C0278818|T191|Recurrent Adrenocortical Carcinoma
C0278818|T191|Recurrent Adrenal Cortex Cancer
C0278818|T191|recurrent adrenocortical carcinoma
C0278818|T191|Relapsed Carcinoma of Adrenal Cortex
C0278818|T191|Recurrent Carcinoma of Adrenal Cortex
C0278818|T191|recurrent adrenocortical cancer
C0278818|T191|Relapsed Adrenal Cortex Carcinoma
C0278818|T191|carcinoma, adrenocortical recurrent
C1709929|T049|Restriction Site Polymorphism
C1881237|T061|Interstitial Radiation Therapy
C1881237|T061|interstitial radiation therapy
C1881237|T061|implant radiation
C1881237|T061|Implant Radiation
C2985558|T061|High-energy Photon Therapy
C2985558|T061|high-energy photon therapy
CL448399|T191|Recurrent Urothelial Carcinoma of the Renal Pelvis and Ureter
CL448399|T191|Relapsed Transitional Cell Cancer of Renal Pelvis and Ureter
CL448399|T191|Relapsed Transitional Cell Carcinoma of the Renal Pelvis and Ureter
CL448399|T191|Relapsed Transitional Cell Cancer of the Renal Pelvis and Ureter
CL448399|T191|Recurrent Transitional Cell Cancer of the Renal Pelvis and Ureter
CL448399|T191|Relapsed Transitional Cell Carcinoma of Renal Pelvis and Ureter
CL448399|T191|Recurrent Transitional Cell Cancer of Renal Pelvis and Ureter
CL448399|T191|Recurrent Transitional Cell Carcinoma of Renal Pelvis and Ureter
C1514422|T191|Primary Glioblastoma
C1514422|T191|Primary Glioblastoma Multiforme
C1517894|T191|Lipid-Rich Breast Carcinoma
C1517894|T191|Lipid Secreting Breast Carcinoma
C0855096|T191|Recurrent Small Lymphocytic Lymphoma
C0855096|T191|Relapsed B-Cell Small Lymphocytic Lymphoma
C0855096|T191|B-cell small lymphocytic lymphoma recurrent
C0855096|T191|Small lymphocyte B lymphoma (Lukes-Collins Classification) recurrent
C0855096|T191|Relapsed Small Lymphocytic Lymphoma
C0855096|T191|Recurrent B-Cell Small Lymphocytic Lymphoma
C0855096|T191|small lymphocytic lymphoma, relapsed
C0855096|T191|recurrent small lymphocytic lymphoma
C0855096|T191|small lymphocytic lymphoma, recurrent
C0855096|T191|relapsed small lymphocytic lymphoma
C106076|T061|Tandem Brachytherapy
C0404187|T061|Left Salpingo-Oophorectomy
C1519323|T049|Silent Mutation
C1519323|T049|Exonic Synonymous Mutation
C1519323|T049|Mutation, Silent
C1519323|T049|Exon Synonymous Mutation
C1519323|T049|Synonymous Mutation
C0149614|T190|Adnexal Mass
C0149614|T190|adnexal mass
C0149614|T190|Adnexal mass
C0149614|T190|ADNEXAL MASS
C1514471|T034|Progesterone Receptor Status
C1514471|T034|PgR Status
C030852|T121|Vinorelbine
C030852|T121|nor-5'-Anhydrovinblastine
C030852|T121|3',4'-Didehydro-4'-deoxy-C'-norvincaleukoblastine
C030852|T121|VNB
C030852|T121|Dihydroxydeoxynorvinkaleukoblastine
C030852|T121|NVB
C030852|T121|Vinorelbine (substance)
C030852|T121|Eunades
C030852|T121|608210
C030852|T121|Biovelbin
C030852|T121|vinorelbine [Chemical/Ingredient]
C030852|T121|navelbine ditartrate
C030852|T121|5'-Nor-Anhydrovinblastine
C030852|T121|C'-Norvincaleukoblastine, 3',4'-didehydro-4'-deoxy-
C030852|T121|vinorelbine
C030852|T121|5'-nor-anhydrovinblastine
C030852|T121|VINORELBINE
C030852|T121|Vinorelbine (product)
C0278554|T191|Recurrent Rectal Carcinoma
C0278554|T191|Rectal carcinoma recurrent
C0278554|T191|recurrent rectal cancer
C0278554|T191|Rectal cancer recurrent
C0278554|T191|Recurrent Cancer of Rectum
C0278554|T191|Carcinoma rectum recurrent
C0278554|T191|rectal cancer, recurrent
C0278554|T191|Recurrent Rectal Cancer
C0278554|T191|Recurrent Cancer of the Rectum
C0278554|T191|Rectal Cancer, Recurrent
C0278554|T191|rectum cancer, recurrent
C0278554|T191|Carcinoma of rectum recurrent
C0278554|T191|recurrent rectum cancer
C3273215|T191|Invasive Lobular Breast Carcinoma, Alveolar Variant
C1332347|T191|Atypical Ductal Breast Hyperplasia
C1332347|T191|Atypical hyperplasia of lactiferous duct (disorder)
C1332347|T191|Ductal Intraepithelial Neoplasia, Grade 1B
C1332347|T191|Atypical ductal hyperplasia of breast
C1332347|T191|Atypical Ductal Hyperplasia of Breast
C1332347|T191|Atypical Breast Ductal Hyperplasia
C1332347|T191|ADH
C1332347|T191|Atypical mammary duct hyperplasia
C1332347|T191|DIN 1B
C1332347|T191|Atypical hyperplasia of lactiferous duct
C1332347|T191|atypical ductal breast hyperplasia
C1332347|T191|atypical ductal hyperplasia
C1332347|T191|Atypical Ductal Hyperplasia of the Breast
C1514512|T191|Prostate Ductal Adenocarcinoma, Papillary Pattern
C0278680|T191|Localized Parathyroid Gland Carcinoma
C0278680|T191|parathyroid cancer, localized
C0278680|T191|carcinoma of the parathyroid, localized
C0278680|T191|parathyroid carcinoma, localized
C0278680|T191|localized parathyroid cancer
C0278680|T191|localized parathyroid carcinoma
C0278680|T191|Localized Parathyroid Carcinoma
C0278680|T191|cancer of the parathyroid, localized
C0278680|T191|Localized Parathyroid Cancer
C1336882|T191|Infiltrating Ureter Urothelial Carcinoma with Squamous Differentiation
C1336882|T191|Transitional Cell Carcinoma of Ureter with Squamous Differentiation
C1336882|T191|Transitional Cell Carcinoma of the Ureter with Squamous Differentiation
C1336882|T191|Ureteral Transitional Cell Carcinoma with Squamous Differentiation
C1881249|T045|Intron Splice Region Mutation
C1881249|T045|Splice Region Mutation
C1881249|T045|Intronic Splice Region Mutation
C1335661|T191|Radiation-Related Angiosarcoma
C1335661|T191|Radiation-Induced Angiosarcoma
C1332998|T191|Childhood T Lymphoblastic Lymphoma
C1332998|T191|Childhood Precursor T-Lymphoblastic Lymphoma
C0686617|T191|Metastatic Malignant Neoplasm to the Thymus
C0686617|T191|Metastatic Tumor to the Thymus
C0686617|T191|Secondary Malignant Tumor to the Thymus
C0686617|T191|Metastatic Neoplasm to the Thymus
C0686617|T191|Metastatic Malignant Tumor to the Thymus
C0686617|T191|Metastasis to the Thymus
C0686617|T191|Secondary Malignant Neoplasm to the Thymus
C1514506|T191|Prostate Adenocarcinoma with Focal Neuroendocrine Differentiation
C0278776|T191|Recurrent Childhood Acute Myeloid Leukemia
C0278776|T191|relapsed pediatric acute nonlymphocytic leukemia
C0278776|T191|childhood acute myeloid leukemia, relapsed
C0278776|T191|Recurrent Childhood Acute Myelocytic Leukemia
C0278776|T191|acute myeloid leukemia, relapsed, childhood
C0278776|T191|childhood AML, relapsed
C0278776|T191|Relapsed Pediatric Acute Myelogenous Leukemia
C0278776|T191|recurent childhood AML
C0278776|T191|Relapsed Childhood Acute Myeloblastic Leukemia
C0278776|T191|recurrent pediatric acute myeloid leukemia
C0278776|T191|leukemia, recurrent childhood acute myeloid
C0278776|T191|childhood leukemia, acute nonlymphocytic relapsed
C0278776|T191|Recurrent Childhood Acute Myeloblastic Leukemia
C0278776|T191|pediatric leukemia, acute myeloid relapsed
C0278776|T191|acute nonlymphocytic leukemia, relapsed, childhood
C0278776|T191|Recurrent Pediatric Acute Myeloblastic Leukemia
C0278776|T191|myeloid leukemia, relapsed childhood acute
C0278776|T191|recurrent childhood ANLL
C0278776|T191|childhood AML, recurrent
C0278776|T191|pediatric acute myeloid leukemia, relapsed
C0278776|T191|Relapsed Childhood Acute Myelogenous Leukemia
C0278776|T191|Relapsed Pediatric Acute Myeloid Leukemia
C0278776|T191|recurrent childhood acute nonlymphocytic leukemia
C0278776|T191|nonlymphocytic leukemia, relapsed pediatric acute
C0278776|T191|leukemia, reucrrent childhood acute nonlymphocytic
C0278776|T191|childhood acute nonlymphocytic leukemia, relapsed
C0278776|T191|nonlymphocytic leukemia, relapsed childhood acute
C0278776|T191|Recurrent Pediatric Acute Myelocytic Leukemia
C0278776|T191|relapsed childhood AML
C0278776|T191|Recurrent Childhood Acute Myelogenous Leukemia
C0278776|T191|relapsed childhood acute myeloid leukemia
C0278776|T191|Recurrent Pediatric AML
C0278776|T191|ANLL, recurrent, pediatric
C0278776|T191|AML, recurrent, childhood
C0278776|T191|relapsed pediatric acute myeloid leukemia
C0278776|T191|AML, relapsed, pediatric
C0278776|T191|acute myeloid leukemia, recurrent, childhood
C0278776|T191|pediatric leukemia, acute nonlymphocytic relapsed
C0278776|T191|Relapsed Pediatric Acute Myeloblastic Leukemia
C0278776|T191|Relapsed Childhood Acute Myeloid Leukemia
C0278776|T191|Recurrent Childhood AML
C0278776|T191|relapsed childhood ANLL
C0278776|T191|relapsed pediatric ANLL
C0278776|T191|myeloid leukemia, relapsed pediatric acute
C0278776|T191|ANLL, relapsed, pediatric
C0278776|T191|recurrent pediatric acute nonlymphocytic leukemia
C0278776|T191|Recurrent Pediatric Acute Myeloid Leukemia
C0278776|T191|Relapsed Pediatric AML
C0278776|T191|recurrent childhood acute myeloid leukemia
C0278776|T191|childhood acute myeloid leukemia, recurrent
C0278776|T191|Relapsed Childhood AML
C0278776|T191|Recurrent Pediatric Acute Myelogenous Leukemia
C0278776|T191|Relapsed Childhood Acute Myelocytic Leukemia
C0278776|T191|Recurrent Childhood Acute Non-Lymphocytic Leukemia
C0278776|T191|relapsed pediatric AML
C0278776|T191|relapsed childhood acute nonlymphocytic leukemia
C0278776|T191|AML, relapsed, childhood
C0278776|T191|leukemia, relapsed childhood acute nonlymphocytic
C0278776|T191|ANLL, relapsed, childhood
C0278776|T191|ANLL, recurrent, childhood
C0278776|T191|Relapsed Pediatric Acute Myelocytic Leukemia
C0278776|T191|childhood leukemia, acute myeloid relapsed
C0278776|T191|AML, recurrent, pediatric
C0278776|T191|pediatric acute nonlymphocytic leukemia, relapsed
C0278776|T191|leukemia, relapsed childhood acute myeloid
C0855053|T191|Recurrent Extraskeletal Osteosarcoma
C0855053|T191|Recurrent Extraosseous Osteosarcoma
C0855053|T191|Recurrent Extraskeletal Osteogenic Sarcoma
C0855053|T191|Relapsed Extraskeletal Osteosarcoma
C0855053|T191|Extraskeletal Osteosarcoma, Recurrent
C0855053|T191|Relapsed Extraskeletal Osteogenic Sarcoma
C0855053|T191|Extraskeletal osteosarcoma recurrent
C0262613|T033|Renal Mass
C0262613|T033|Kidney Mass
C0262613|T033|Renal mass NOS
C0262613|T033|KIDNEY MASS
C0262613|T033|Kidney mass
C0262613|T033|Renal mass (finding)
C0262613|T033|Renal mass
C0262613|T033|RENAL MASS
C0347003|T191|Metastatic Malignant Neoplasm to the Testis
C0347003|T191|Metastatic Tumor to the Testis
C0347003|T191|Metastatic Neoplasm to the Testis
C1332234|T191|Alkylating Agent-Related Acute Myeloid Leukemia and Myelodysplastic Syndrome
C1332234|T191|Alkylating Agent-Related AML and MDS
C1332234|T191|Alkylating Agent Related Acute Myeloid Leukemia and Myelodysplastic Syndrome
C0290883|T121|Anastrozole
C0290883|T121|Alpha,alpha,alpha', alpha'-tetramethyl-5-(1H-1,2,4-triazol-1-ylmethyl)-1,3-benzenediacetonitrile
C0290883|T121|2,2'-[5-(1H-1,2,4-Triazol-1-ylmethyl)-1,3-phenylene]di(2-methylpropionitrile)
C0290883|T121|ZD-1033
C0290883|T121|ICI-D1033
C0290883|T121|ANASTROZOLE
C0290883|T121|Arimidex
C0290883|T121|anastrozole
C0290883|T121|ICI D1033
C0347016|T191|Metastatic Malignant Neoplasm to the Spinal Cord
C0347016|T191|Metastatic Neoplasm to the Spinal Cord
C0347016|T191|Metastasis to Spinal Cord
C0347016|T191|Secondary Malignant Neoplasm to the Spinal Cord
C0347016|T191|Metastatic Tumor to the Spinal Cord
C0347016|T191|Secondary Malignant Tumor to the Spinal Cord
C1334708|T191|Metaplastic Breast Carcinoma
C1334708|T191|Metaplastic Carcinoma of Breast
C1334708|T191|Metaplastic breast carcinoma
C1334708|T191|Metaplastic Carcinoma of the Breast
C1334274|T191|Invasive Carcinoma
C2698750|T191|Pediatric Follicular Lymphoma
C2698750|T191|Childhood Follicular Lymphoma
C0010583|T121|Cyclophosphamide
C0010583|T121|CPM - cyclophosphamide
C0010583|T121|N,N-bis(2-chloroethyl)-N',O-propylenephosphoric acid ester diamide monohydrate
C0010583|T121|Genoxal
C0010583|T121|Cytophosphane
C0010583|T121|N,N-bis(beta-chloroethyl)-N',O-propylenephosphoric acid ester diamide monohydrate
C0010583|T121|Endoxana
C0010583|T121|Cyclophosphamidum
C0010583|T121|4173
C0010583|T121|cyclophosphamide
C0010583|T121|Sendoxan
C0010583|T121|Bis(2-chloroethyl)phosphoramide cyclic propanolamide ester monohydrate
C0010583|T121|N,N-bis(2-chloroethyl)tetrahydro-2H-1,3,2-oxazaphosphorin-2-amine 2-oxide monohydrate
C0010583|T121|2-[bis(2-chloroethyl)amino]tetrahydro-2H-1,3,2-oxazaphosphorine 2-oxide monohydrate
C0010583|T121|Cytophosphan
C0010583|T121|CPM
C0010583|T121|Fosfaseron
C0010583|T121|Enduxan
C0010583|T121|B-518
C0010583|T121|(-)-Cyclophosphamide
C0010583|T121|Mitoxan
C0010583|T121|Ciclofosfamida
C0010583|T121|Neosar
C0010583|T121|2-[bis(b-chloroethyl)amino]-1-oxa-3-aza-2-phosphacyclohexane-2-oxide monohydrate
C0010583|T121|Monohydrate, Cyclophosphamide
C0010583|T121|Procytox
C0010583|T121|CP monohydrate
C0010583|T121|CYT
C0010583|T121|Cyclostine
C0010583|T121|Cyclophosphamid monohydrate
C0010583|T121|6055-19-2 (monohydrate)
C0010583|T121|Endoxan
C0010583|T121|Cyclophosphamide (substance)
C0010583|T121|7089
C0010583|T121|Ledoxina
C0010583|T121|Genuxal
C0010583|T121|Cycloblastin
C0010583|T121|bis(2-chloroethyl)phosphamide cyclic propanolamide ester monohydrate
C0010583|T121|N,N-bis(b-chloroethyl)-N',O-trimethylenephosphoric acid ester diamide monohydrate
C0010583|T121|Cyclostin
C0010583|T121|26271
C0010583|T121|Zytoxan
C0010583|T121|WR-138719
C0010583|T121|Cyclophosphamide [Chemical/Ingredient]
C0010583|T121|Cycloblastine
C0010583|T121|Cytoxan
C0010583|T121|Cyclophospham
C0010583|T121|Cyclophosphane
C0010583|T121|Carloxan
C0010583|T121|CYCLO-cell
C0010583|T121|Cicloxal
C0010583|T121|2-[di(chloroethyl)amino]-1-oxa-3-aza-2-phosphacyclohexane 2-oxide monohydrate
C0010583|T121|2H-1,3,2-Oxazaphosphorin-2-amine, N,N-bis(2-chloroethyl)tetrahydro-, 2-oxide
C0010583|T121|CYCLOPHOSPHAMIDE
C0010583|T121|Cyclophosphamide Monohydrate
C0010583|T121|2H-1,3,2-Oxazaphosphorine, 2-[bis(2-chloroethyl)amino]tetrahydro-, 2-oxide, monohydrate
C0010583|T121|1-bis(2-chloroethyl)-amino-1-oxo-2-aza-5-oxaphosphoridin monohydrate
C0010583|T121|Clafen
C0010583|T121|CTX
C0010583|T121|bis(2-chloroethyl)phosphoramide cyclic propanolamide ester monohydrate
C0010583|T121|Ciclofosfamide
C0010583|T121|N,N-bis(2-chloroethyl)-N'-(3-hydroxypropyl)phosphorodiamidic acid intramolecular ester monohydrate
C0010583|T121|CTX - cyclophosphamide
C0010583|T121|N,N-bis(beta-chloroethyl)-N',O-trimethylenephosphoric acid ester diamide monohydrate
C0010583|T121|Cyclophosphanum
C0010583|T121|Cyclophosphan
C0010583|T121|Cyclophosphamide (product)
C0010583|T121|Asta B 518
C0010583|T121|CYT - cyclophosphamide
C0010583|T121|WR- 138719
C0010583|T121|Claphene
C0010583|T121|Syklofosfamid
C1336536|T191|Supratentorial Glioblastoma
C1336536|T191|Supratentorial Glioblastoma Multiforme
C1336536|T191|Grade IV Supratentorial Astrocytic Tumor
C1336536|T191|Grade IV Supratentorial Astrocytic Neoplasm
C1334417|T191|Low Grade Mucoepidermoid Breast Carcinoma
C1334417|T191|Low-Grade Mucoepidermoid Carcinoma of the Breast
C1334417|T191|Low-Grade Mucoepidermoid Carcinoma of Breast
C0039286|T121|Tamoxifen
C0039286|T121|Ethanamine, 2-(4-(1,2-diphenyl-1-butenyl)phenoxy)-N,N-dimethyl-, (Z)-
C0039286|T121|TAMOXIFEN
C0039286|T121|TAM
C0039286|T121|(Z)-2-[4-(1,2-diphenyl-1-butenyl)phenoxy]-N,N-dimethylethanamine 2-hydroxy-1,2,3-propanetricarboxylate (1:1)
C0039286|T121|Tamoxifen [Chemical/Ingredient]
C0039286|T121|tamoxifen
C0039286|T121|TMX
C0039286|T121|Tamoxifen (product)
C0039286|T121|1-p-beta-dimethylamino-ethoxyphenyl-trans-1,2-diphenylbut-1-ene
C0039286|T121|Tamoxifen (substance)
C0728747|T116|Trastuzumab
C0728747|T116|Anti-erbB-2
C0728747|T116|Monoclonal Antibody c-erb-2
C0728747|T116|MoAb HER2
C0728747|T116|Anti-p185-HER2
C0728747|T116|c-erb-2 Monoclonal Antibody
C0728747|T116|Herceptin Biosimilar PF-05280014
C0728747|T116|Anti-erbB2 Monoclonal Antibody
C0728747|T116|Anti-ERB-2
C0728747|T116|Herceptin Trastuzumab Biosimilar PF-05280014
C0728747|T116|Trastuzumab Biosimilar ABP 980
C0728747|T116|TRASTUZUMAB
C0728747|T116|trastuzumab
C0728747|T116|ABP 980
C0728747|T116|PF-05280014
C0728747|T116|Trastuzumab Biosimilar PF-05280014
C0728747|T116|Anti-c-ERB-2
C0728747|T116|Anti-c-erbB2 Monoclonal Antibody
C0728747|T116|rhuMAb HER2
C0728747|T116|Anti-HER2/c-erbB2 Monoclonal Antibody
C0728747|T116|HER2 Monoclonal Antibody
C0728747|T116|Monoclonal Antibody HER2
C0728747|T116|Herceptin
C0853826|T191|Anaplastic (Malignant) Intraspinal Meningioma
C0853826|T191|Malignant Meningioma of Spinal Canal and Spinal Cord
C0853826|T191|Malignant Intraspinal Meningioma
C0853826|T191|Malignant Spinal Canal and Spinal Cord Meningioma
C0853826|T191|Malignant Meningioma of the Spinal Canal and Spinal Cord
C0853826|T191|Anaplastic Intraspinal Meningioma
C2945703|T061|Prophylactic Oophorectomy
C2945703|T061|prophylactic oophorectomy
C0475385|T185|T1b Stage Finding
C0475385|T185|T1b Primary Tumor Stage Finding
C0475385|T185|T1b
C0475385|T185|Tumor stage T1b
C0475385|T185|T1b Stage
C0475385|T185|T1b Primary Tumor Finding
C0475385|T185|T1b TNM Finding
C0475385|T185|T1b Tumor Finding
C0475385|T185|Tumor Stage T1b
C0475385|T185|Tumor stage T1b (finding)
C0475385|T185|T1b Cancer Stage Finding
C0475385|T185|T1b Tumor Stage
C0475385|T185|Tumour stage T1b
C1266043|T191|Sarcomatoid Renal Cell Carcinoma
C1266043|T191|RCC w/ sarcomatoid features
C1266043|T191|Renal cell carcinoma, sarcomatoid
C1266043|T191|Renal cell carcinoma, spindle cell
C1266043|T191|Renal cell carcinoma, sarcomatoid (morphologic abnormality)
C1266043|T191|Renal cell carcinoma with sarcomatoid features
C0853709|T191|Recurrent Lymphoplasmacytic Lymphoma
C0853709|T191|Lymphoplasmacytoid immunocytoma recurrent
C0853709|T191|Lymphoplasmacytoid lymphoma/immunocytoma recurrent
C0853709|T191|Waldenstrom's macroglobulinemia recurrent
C0853709|T191|Relapsed Lymphoplasmacytoid Lymphoma/Immunocytoma
C0853709|T191|Immunocytoma (Lymphoplasmacytoid lymphoma/immunocytoma) (Kiel Classification) recurrent
C0853709|T191|Recurrent Lymphoplasmacytoid Lymphoma/Immunocytoma
C0853709|T191|Waldenstrom's macroglobulinaemia recurrent
C0855069|T191|Recurrent Rhabdomyosarcoma
C0855069|T191|Rhabdosarcoma recurrent
C0855069|T191|Relapsed Rhabdomyosarcoma
C0855069|T191|Rhabdomyosarcoma Recurrent
C0855069|T191|Rhabdomyosarcoma recurrent
C0280190|T191|Recurrent Adult Immunoblastic Lymphoma
C0280190|T191|Recurrent Adult Immunoblastic Large Cell Lymphoma
C0280190|T191|immunoblastic large cell lymphoma, recurrent, adult
C0280190|T191|adult immunoblastic large cell lymphoma, recurrent
C0280190|T191|Relapsed Adult Immunoblastic Lymphoma
C0280190|T191|adult immunoblastic large cell lymphoma, relapsed
C0280190|T191|recurrent adult immunoblastic large cell lymphoma
C0280190|T191|relapsed adult immunoblastic large cell lymphoma
C0280190|T191|immunoblastic large cell lymphoma, adult, recurrent
C0280190|T191|Relapsed Adult Immunoblastic Large Cell Lymphoma
C2350866|T121|Eribulin
C2350866|T121|ER-086526
C2350866|T121|2-(3-amino-2-hydroxypropyl)hexacosahydro-3-methoxy-26-methyl-20,27-bis(methylene)11,15-18,21-24,28-triepoxy-7,9-ethano-12,15-methano-9H,15H-furo(3,2-i)furo(2',3'-5,6)pyrano(4,3-b)(1,4)dioxacyclopentacosin-5-(4H)-one
C2350866|T121|2-(3-Amino-2-hydroxypropyl)hexacosahydro-3-methoxy-26-methyl-20,27-bis(methylene)11,15-18,21-24,28-triepoxy-7,9-ethano-12,15-methano-9H,15H-furo(3,2-i)furo(2',3'-5,6)pyrano(4,3-b)(1,4)dioxacyclopentacosin-5-(4H)-one
C2350866|T121|ERIBULIN
C2350866|T121|eribulin
C0278739|T191|Recurrent Childhood Lymphoblastic Lymphoma
C0278739|T191|Relapsed Childhood Lymphoblastic Lymphoma
C0278739|T191|recurrent lymphoblastic childhood lymphoma
C0278739|T191|lymphoma, non-Hodgkin's, lymphoblastic recurrent, childhood
C0278739|T191|non-Hodgkin's lymphoma, lymphoblastic recurrent, childhood
C0278739|T191|Recurrent Pediatric Lymphoblastic Lymphoma
C0278739|T191|pediatric lymphoblastic non-Hodgkin's lymphoma, recurrent
C0278739|T191|childhood non-Hodgkin's lymphoma, lymphoblastic recurrent
C0278739|T191|lymphoblastic recurrent non-Hodgkin's lymphoma, childhood
C0278739|T191|relapsed lymphoblastic childhood lymphoma
C0278739|T191|relapsed childhood lymphoblastic lymphoma
C0278739|T191|Relapsed Pediatric Lymphoblastic Lymphoma
C0278739|T191|Recurrent Childhood Precursor Lymphoblastic Lymphoma
C0278739|T191|NHL, lymphoblastic recurrent childhood
C0278739|T191|recurrent childhood lymphoblastic lymphoma
C0862417|T191|Stage III Bladder Urothelial Carcinoma
C0862417|T191|Stage III Transitional Cell Carcinoma of Bladder
C0862417|T191|Stage III Transitional Cell Carcinoma of the Bladder
C0862417|T191|Stage III Bladder Urothelial Carcinoma AJCC v6
C0862417|T191|Stage III Transitional Cell Carcinoma of the Urinary Bladder
C0862417|T191|Stage III Bladder Urothelial Carcinoma AJCC v7
C0862417|T191|Stage III Urinary Bladder Transitional Cell Carcinoma
C0862417|T191|Stage III Transitional Cell Carcinoma of Urinary Bladder
C1708718|T191|Localized Non-Resectable Adult Hepatocellular Carcinoma
C1708718|T191|Localized Unresectable Adult Hepatocellular Carcinoma
C1300499|T201|Tumor size, dominant nodule, greatest dimension, in specimen obtained by prostatic enucleation
C1300499|T201|Tumour size, dominant nodule, greatest dimension, in specimen obtained by prostatic enucleation
C1300499|T201|Tumor size, dominant nodule, greatest dimension, in specimen obtained by prostatic enucleation (observable entity)
C1515024|T191|Submucosal Invasive Colon Adenocarcinoma
C1706716|T049|Adenosine to Cytosine Transversion Abnormality
C1706716|T049|Adenosine to Cytosine Mutation
C1706716|T049|Adenosine to Cytosine Transversion
C0041692|T061|Unilateral Salpingo-oophorectomy
C0041692|T061|unilateral salpingo-oophorectomy
C0334588|T191|Giant Cell Glioblastoma
C0334588|T191|Giant Cell Glioblastomas
C0334588|T191|Giant cell glioblastoma (morphologic abnormality)
C0334588|T191|giant cell glioblastoma (WHO grade IV)
C0334588|T191|Giant cell glioblastoma
C0334588|T191|giant cell glioblastoma
C0334588|T191|Glioblastoma, Giant Cell
C0334588|T191|Monstrocellular sarcoma [obs]
C0334588|T191|Glioblastomas, Giant Cell
C0854866|T191|Recurrent Non-Hodgkin Lymphoma
C0854866|T191|Relapsed Non-Hodgkin's Lymphoma
C0854866|T191|Non-Hodgkin's Lymphoma Relapsed
C0854866|T191|Recurrent Non-Hodgkin's Lymphoma
C0854761|T191|Recurrent Esophageal Carcinoma
C0854761|T191|Relapsed Carcinoma of Esophagus
C0854761|T191|Recurrent Carcinoma of the Esophagus
C0854761|T191|Recurrent Cancer of the Esophagus
C0854761|T191|Relapsed Esophageal Cancer
C0854761|T191|Esophageal Carcinoma, Recurrent
C0854761|T191|Relapsed Cancer of the Esophagus
C0854761|T191|Recurrent Esophageal Cancer
C0854761|T191|Relapsed Esophagus Carcinoma
C0854761|T191|Recurrent Cancer of Esophagus
C0854761|T191|Recurrent Carcinoma of Esophagus
C0854761|T191|Oesophageal carcinoma site unspecified recurrent
C0854761|T191|Oesophageal carcinoma recurrent
C0854761|T191|Esophageal carcinoma site unspecified recurrent
C0854761|T191|esophagus cancer, recurrent
C0854761|T191|Relapsed Cancer of Esophagus
C0854761|T191|recurrent esophageal cancer
C0854761|T191|Esophageal carcinoma recurrent
C0854761|T191|esophageal cancer, recurrent
C0854761|T191|Oesophageal Carcinoma Recurrent
C0854761|T191|Relapsed Carcinoma of the Esophagus
C0854761|T191|Recurrent Esophagus Cancer
C0279087|T191|Recurrent Kaposi Sarcoma
C0279087|T191|Kaposi's sarcoma, recurrent
C0279087|T191|sarcoma, multiple hemorrhagic, recurrent
C0279087|T191|Recurrent Kaposi's Sarcoma
C0279087|T191|multiple hemorrhagic sarcoma, recurrent
C0279087|T191|recurrent multiple hemorrhagic sarcoma
C0279087|T191|recurrent Kaposi sarcoma
C0279087|T191|Recurrent Multiple Hemorrhagic Sarcoma
C0279087|T191|sarcoma, Kaposi's, recurrent
C0441916|T033|LX stage
C0441916|T033|LX
C0441916|T033|LX Stage
C0441916|T033|Lymphatic Stage LX
C0441916|T033|Lymphatic stage LX
C0441916|T033|LX TNM Finding
C0441916|T033|LX Lymphatic Vessel Invasion Finding
C0441916|T033|LX Lymphatic Stage
C0441916|T033|LX: lymphatic vessel invasion cannot be assessed
C0441916|T033|LX Lymphatic Invasion Finding
C0441916|T033|LX Stage Finding
C0441916|T033|LX Cancer Stage Finding
C0441916|T033|LX stage (finding)
C1883645|T086|5' Untranslated Region Mutation
C1883645|T086|5' UTR Mutation
CL412336|T061|Microwave Ablation
CL412336|T061|microwave ablation
C1306459|T191|Primary Malignant Neoplasm
C1306459|T191|Malignant neoplasm, primary (morphologic abnormality)
C1306459|T191|Blastoma
C1306459|T191|Malignant neoplasm
C1306459|T191|Malignant tumor morphology
C1306459|T191|Neoplasm, malignant
C1306459|T191|Primary malignant neoplasm (disorder)
C1306459|T191|Cancer
C1306459|T191|Unclassified tumour, malignant
C1306459|T191|Tumor, malignant
C1306459|T191|Tumour, malignant
C1306459|T191|Malignancy
C1306459|T191|Neoplasm, malignant (primary)
C1306459|T191|Cancer morphology
C1306459|T191|Malignant neoplasm, primary
C1306459|T191|Malignant tumour morphology
C1306459|T191|Unclassified tumor, malignant
C1306459|T191|Primary malignant neoplasm
C1708063|T061|First-Line Therapy
C1708063|T061|First-Line Treatment
C1708063|T061|primary treatment
C1708063|T061|First Line Treatment
C1708063|T061|primary therapy
C1708063|T061|First Line Therapy
C1708063|T061|first-line therapy
C1710347|T049|Tandem Repeat Variation
C1710347|T049|VNTR
C1710347|T049|Variable Number Tandem Repeat
C0854638|T061|Antiestrogen Therapy
C0854638|T061|Antiestrogen therapy
C0854638|T061|Antioestrogen therapy
C0854638|T061|antiestrogen therapy
C0854638|T061|therapy, antiestrogen
C0206726|T191|Gliosarcoma
C0206726|T191|Glioblastoma with a Sarcomatous Component
C0206726|T191|Sarcomatous Glioma
C0206726|T191|Gliosarcomas
C0206726|T191|Sarcomatous Gliomas
C0206726|T191|gliosarcoma (WHO grade IV)
C0206726|T191|gliosarcoma
C0206726|T191|Glioma, Sarcomatous
C0206726|T191|Gliosarcoma (morphologic abnormality)
C0206726|T191|Glioblastoma with Sarcomatous Component
C0206726|T191|Gliosarcoma [Disease/Finding]
C0206726|T191|Glioblastoma with sarcomatous component
C0206726|T191|Gliomas, Sarcomatous
C0686507|T191|Metastatic Malignant Neoplasm to the Parathyroid Gland
C0686507|T191|Metastatic Neoplasm to the Parathyroid
C0686507|T191|Metastatic Neoplasm to the Parathyroid Gland
C0686507|T191|Metastatic Tumor to the Parathyroid Gland
C0686507|T191|Metastasis to the Parathyroid Gland
C0686507|T191|Metastatic Tumor to the Parathyroid
C1519214|T191|Secondary Glioblastoma
C1519214|T191|Secondary Glioblastoma Multiforme
C0751366|T191|Radiation-Related Malignant Neoplasm
C0751366|T191|Radiation-Induced Cancer
C0751366|T191|Radiation-Related Cancer
C0751366|T191|Radiation-Induced Malignant Neoplasm
C1880435|T061|EC Breast Regimen
C1880435|T061|Epirubicin-Cytoxan Regimen
C0862490|T191|Metastatic Endometrioid Adenocarcinoma
C0862490|T191|Endometrioid adenocarcinoma metastatic
C0862490|T191|Metastatic Endometrioid Carcinoma
C0279988|T191|Childhood Angiosarcoma
C0279988|T191|Pediatric Hemangiosarcoma
C0279988|T191|hemangiosarcoma, childhood
C0279988|T191|Pediatric Angiosarcoma
C0279988|T191|hemangiosarcoma, pediatric
C0279988|T191|pediatric angiosarcoma
C0279988|T191|sarcoma, angio-, pediatric
C0279988|T191|childhood hemangiosarcoma
C0279988|T191|angiosarcoma, childhood
C0279988|T191|pediatric hemangiosarcoma
C0279988|T191|childhood angiosarcoma
C0279988|T191|angiosarcoma, pediatric
C0279988|T191|sarcoma, angio-, childhood
C0279988|T191|Childhood Hemangiosarcoma
C1334587|T191|Growth Hormone-Producing Pituitary Gland Carcinoma
C1334587|T191|Malignant Somatotropinoma of Pituitary
C1334587|T191|Malignant Growth Hormone Producing Tumor of the Pituitary
C1334587|T191|Malignant Growth Hormone Producing Neoplasm of the Pituitary Gland
C1334587|T191|Malignant Growth Hormone Secreting Neoplasm of the Pituitary
C1334587|T191|Malignant Growth Hormone Secreting Tumor of the Pituitary
C1334587|T191|Malignant Pituitary Gland Somatotropinoma
C1334587|T191|Malignant Growth Hormone Producing Pituitary Gland Tumor
C1334587|T191|Growth Hormone Producing Pituitary Gland Carcinoma
C1334587|T191|Malignant Growth Hormone Secreting Neoplasm of Pituitary Gland
C1334587|T191|Malignant Growth Hormone Secreting Tumor of Pituitary
C1334587|T191|Malignant Pituitary Somatotropinoma
C1334587|T191|Malignant Somatotropinoma of the Pituitary
C1334587|T191|Malignant Growth Hormone Producing Pituitary Neoplasm
C1334587|T191|Malignant Growth Hormone Secreting Pituitary Gland Tumor
C1334587|T191|Malignant Growth Hormone Secreting Tumor of the Pituitary Gland
C1334587|T191|Malignant Growth Hormone Producing Tumor of Pituitary Gland
C1334587|T191|Malignant Somatotropinoma of the Pituitary Gland
C1334587|T191|Malignant Growth Hormone Producing Tumor of the Pituitary Gland
C1334587|T191|Malignant Growth Hormone Producing Neoplasm of Pituitary Gland
C1334587|T191|Malignant Growth Hormone Secreting Pituitary Tumor
C1334587|T191|Malignant Growth Hormone Producing Neoplasm of the Pituitary
C1334587|T191|Malignant Growth Hormone Producing Pituitary Gland Neoplasm
C1334587|T191|Malignant Growth Hormone Secreting Neoplasm of the Pituitary Gland
C1334587|T191|Malignant Growth Hormone Secreting Neoplasm of Pituitary
C1334587|T191|Malignant Growth Hormone Secreting Pituitary Gland Neoplasm
C1334587|T191|Malignant Growth Hormone Producing Neoplasm of Pituitary
C1334587|T191|Malignant Growth Hormone Producing Tumor of Pituitary
C1334587|T191|Malignant Growth Hormone Secreting Tumor of Pituitary Gland
C1334587|T191|Malignant Somatotropinoma of Pituitary Gland
C1334587|T191|Malignant Growth Hormone Producing Pituitary Tumor
C1334587|T191|Malignant Growth Hormone Secreting Pituitary Neoplasm
C1334587|T191|Malignant Growth Hormone Producing Tumor
C2608055|T191|Hereditary Renal Cell Carcinoma
C1883634|T086|3' Untranslated Region Mutation
C1883634|T086|3' UTR Mutation
C1511183|T020|Bistrand Abasic Site
C1333429|T191|Epstein-Barr Virus-Related Clonal Post-Transplant Lymphoproliferative Disorder
C1333429|T191|EBV Related Clonal PTLD
C1333429|T191|EBV-Related Clonal PTLD
C1334716|T191|Metastatic Carcinoma to the Adrenal Cortex
C1334716|T191|Metastatic Carcinoma to Adrenal Cortex
CL448281|T191|Recurrent Nodal Marginal Zone Lymphoma
CL448281|T191|Relapsed Nodal Marginal Zone Lymphoma
CL448281|T191|Recurrent Nodal Marginal Zone B-Cell Lymphoma
C1336924|T191|AIDS-Related Cervical Kaposi Sarcoma
C1336924|T191|AIDS-Related Kaposi's Sarcoma of the Cervix
C1336924|T191|AIDS-Related Cervical Kaposi's Sarcoma
C1336924|T191|AIDS-Related Kaposi's Sarcoma of Cervix
C101267|T034|Estrogen Receptor and/or Progesterone Receptor Positive
C101267|T034|ER and/or PR Positive
C101267|T034|ER and/or PR +
C1882540|T080|Seed Implantation
C1882540|T080|Seed Implant
C1882540|T080|{Seed}
C1882540|T080|Radioactive Seed Implant Dosing Unit
C1882540|T080|Seed
C1882540|T080|radioactive seed
C1882540|T080|seed
C2985437|T049|Null Allele
C2985437|T049|null allele
C1332167|T191|Adenoid Cystic Breast Carcinoma
C1332167|T191|Adenocystic Carcinoma of the Breast
C1332167|T191|Mammary Adenocystic Carcinoma
C1332167|T191|Adenoid cystic breast carcinoma
C1332167|T191|Adenocystic Breast Carcinoma
C1332167|T191|Adenoid Cystic Carcinoma of the Breast
C1332167|T191|Adenoid Cystic Carcinoma of Breast
C1332167|T191|Adenocystic Carcinoma of Breast
C0279647|T191|Childhood Acute Erythroid Leukemia
C0279647|T191|Pediatric Acute Erythroid Leukemia
C0279647|T191|childhood acute M6 leukemia
C0279647|T191|erythroleukemia, childhood acute
C0279647|T191|Pediatric M6 Leukemia
C0279647|T191|pediatric acute erythroleukemia
C0279647|T191|Childhood M6 Leukemia
C0279647|T191|pediatric acute M6 leukemia
C0279647|T191|childhood acute erythroleukemia (M6)
C0279647|T191|leukemia, childhood acute erythro-
C0279647|T191|M6 pediatric acute erythroleukemia
C0279647|T191|M6 leukemia, childhood acute
C0279647|T191|acute erythroleukemia, childhood
C0279647|T191|leukemia, pediatric acute erythro-
C0279647|T191|M6 childhood acute erythroleukemia
C1335737|T191|Recurrent Hematologic Malignancy
C1335737|T191|Relapsed Hematologic Cancer
C1335737|T191|Relapsed Hematologic Malignancy
C1335737|T191|Recurrent Hematologic Cancer
C0346996|T191|Metastatic Malignant Neoplasm to the Cervix
C0346996|T191|Metastasis to the Cervix Uteri
C0346996|T191|Metastasis to the Cervix
C0346996|T191|Metastatic Malignant Tumor to the Uterine Cervix
C0346996|T191|Metastatic Malignant Tumor to the Cervix
C0346996|T191|Metastasis to the Uterine Cervix
C0346996|T191|Metastatic Malignant Neoplasm to the Uterine Cervix
C1333854|T191|Grade 4 Malignant Neoplasm
C0338240|T061|Intraoperative Radiation Therapy
C0338240|T061|radiotherapy, intraoperative
C0338240|T061|IORT
C0338240|T061|Intraoperative radiation therapy
C0338240|T061|Intraoperative Radiotherapy
C0338240|T061|intraoperative radiation therapy
C0338240|T061|intraoperative radiotherapy
C0677798|T061|Thermal Ablation Therapy
C0677798|T061|thermal ablation
C0677798|T061|thermal ablation therapy
C537535|T191|Secretory Breast Carcinoma
C537535|T191|Juvenile Carcinoma of Breast
C537535|T191|Juvenile Secretory Carcinoma of the Breast
C537535|T191|Infiltrating Cystic Hypersecretory Duct Breast Carcinoma
C537535|T191|Secretory breast carcinoma
C537535|T191|Juvenile Secretory Breast Carcinoma
C537535|T191|Invasive Cystic Hypersecretory Duct Breast Carcinoma
C537535|T191|Juvenile Secretory Carcinoma of Breast
C537535|T191|Secretory Carcinoma of the Breast
C537535|T191|Cystic Hypersecretory Carcinoma of the Breast
C537535|T191|Juvenile carcinoma of the breast (morphologic abnormality)
C537535|T191|Secretory Carcinoma of Breast
C537535|T191|Cystic Hypersecretory Breast Carcinoma
C537535|T191|Juvenile Carcinoma of the Breast
C537535|T191|Secretory Carcinoma
C537535|T191|Cystic Hypersecretory Carcinoma of Breast
C537535|T191|Secretory carcinoma of the breast
C537535|T191|Juvenile carcinoma of the breast
C537535|T191|Secretory carcinoma of breast
C537535|T191|Juvenile Breast Carcinoma
C537535|T191|Juvenile carcinoma of breast
C0280674|T061|Aromatase Inhibition Therapy
C0280674|T061|Aromatase inhibition therapy
C0280674|T061|aromatase inhibition therapy
C0280674|T061|inhibition therapy, aromatase
C0280674|T061|Aromatase Inhibition
C1332906|T191|Cerebral Glioblastoma
C1332906|T191|Grade IV Hemispheric Astrocytic Tumor
C1332906|T191|Grade IV Cerebral Hemisphere Astrocytic Tumor
C1332906|T191|Hemispheric Glioblastoma Multiforme
C1332906|T191|Grade IV Astrocytic Tumor of the Cerebral Hemisphere
C1332906|T191|Grade IV Astrocytic Neoplasm of the Cerebral Hemisphere
C1332906|T191|Cerebral Glioblastoma Multiforme
C1332906|T191|Glioblastoma Multiforme of Cerebral Hemisphere
C1332906|T191|Grade IV Astrocytic Neoplasm of Cerebral Hemisphere
C1332906|T191|Glioblastoma Multiforme of the Cerebral Hemisphere
C1332906|T191|Cerebral Hemisphere Glioblastoma Multiforme
C1332906|T191|Grade IV Cerebral Hemisphere Astrocytic Neoplasm
C1332906|T191|Grade IV Hemispheric Astrocytic Neoplasm
C1332906|T191|Grade IV Astrocytic Tumor of Cerebral Hemisphere
CL472691|T191|Childhood Cerebral Anaplastic Astrocytoma
C1300502|T201|Tumor size, dominant nodule, in specimen obtained by radical prostatectomy
C1300502|T201|Tumour size, dominant nodule, in specimen obtained by radical prostatectomy
C1300502|T201|Tumor size, dominant nodule, in specimen obtained by radical prostatectomy (observable entity)
C1520143|T201|Whole-Brain Radiotherapy
C1520143|T201|whole-brain radiation therapy
C1520143|T201|WBRT
C1520143|T201|whole-brain radiotherapy
C1332974|T191|Childhood Conventional Osteosarcoma
C1332974|T191|Childhood Intracortical Osteosarcoma
C1334281|T191|Infiltrating Bladder Urothelial Carcinoma
C1334281|T191|Invasive Bladder Urothelial Carcinoma
C1334281|T191|Infiltrating Transitional Cell Carcinoma of the Urinary Bladder
C1334281|T191|Invasive Transitional Cell Carcinoma of the Urinary Bladder
C1334281|T191|Invasive Bladder Transitional Cell Carcinoma
C1704323|T191|Paget Disease of the Nipple
C1704323|T191|Nipple Paget's Disease
C1704323|T191|Paget's Disease of the Nipple
C1704323|T191|Paget's disease of the nipple
C1704323|T191|Paget's Disease of Nipple
C1882296|T033|Partially Encapsulated Mass
C0861832|T191|Recurrent Duodenal Carcinoma
C0861832|T191|Duodenal carcinoma recurrent
C0861832|T191|Recurrent Duodenal Cancer
C0861832|T191|Duodenal cancer recurrent
C0347020|T191|Metastatic Malignant Neoplasm to the Orbit
C0347020|T191|Metastatic Neoplasm to the Orbit
C0347020|T191|Metastatic Tumor to the Orbit
C0347020|T191|Metastasis to the Orbit
CL376205|T191|Stage IV Childhood Anaplastic Large Cell Lymphoma
CL372028|T191|Childhood Atypical Teratoid/Rhabdoid Tumor
C1334713|T191|Metastatic Bone Ewing Sarcoma
C1334713|T191|Metastatic Ewing's Sarcoma of Bone
C1334713|T191|Metastatic Ewing's Sarcoma of the Bone
C1334713|T191|Metastatic Skeletal Ewing's Sarcoma
C1334713|T191|Metastatic Osseous Ewing's Sarcoma
C1334713|T191|Metastatic Bone Ewing's Sarcoma
C1881801|T191|Metastatic Signet Ring Cell Carcinoma
C1881801|T191|Metastatic signet ring cell carcinoma (morphologic abnormality)
C1881801|T191|Metastatic signet ring cell carcinoma
C1705687|T049|Inversion Mutation Abnormality
C1705687|T049|Inversion Mutation
C1705687|T049|Inversion
C0456906|T033|N1a Stage Finding
C0456906|T033|N1a Regional Lymph Node Stage Finding
C0456906|T033|N1a Lymph Node Finding
C0456906|T033|N1a Regional Lymph Nodes Finding
C0456906|T033|N1a Node Finding
C0456906|T033|Node stage N1a (finding)
C0456906|T033|N1a Cancer Stage Finding
C0456906|T033|N1a TNM Finding
C0456906|T033|N1a Node Stage
C0456906|T033|Lymph Node Stage N1a
C0456906|T033|N1a Stage
C0456906|T033|N1a
C0456906|T033|Node Stage N1a
C0456906|T033|N1a Lymph Node Stage
C0456906|T033|Node stage N1a
C0877373|T191|Advanced Malignant Neoplasm
C0877373|T191|Advanced cancer
C0877373|T191|Advanced Cancer
C0877373|T191|advanced cancer
C1332556|T191|Biphasic Pulmonary Blastoma
C1332556|T191|Classic Pulmonary Blastoma
CL438301|T191|Hereditary Prostate Carcinoma
C0149726|T033|Pulmonary Mass
C0149726|T033|mass
C0149726|T033|Lung mass (finding)
C0149726|T033|Lung Mass
C0149726|T033|Lung mass
C0149726|T033|Pulmonary mass
C0149726|T033|LUNG MASS
C0149726|T033|lung mass
C0347004|T191|Metastatic Malignant Neoplasm to the Epididymis
C0347004|T191|Metastatic Tumor to the Epididymis
C0347004|T191|Metastatic Neoplasm to the Epididymis
C0854977|T191|Recurrent Large Cell Lung Carcinoma
C0854977|T191|Large cell lung cancer recurrent
C0854977|T191|Recurrent Large Cell Carcinoma of the Lung
C0854977|T191|Relapsed Large Cell Lung Carcinoma
C0854977|T191|Recurrent Large Cell Carcinoma of Lung
C0854977|T191|Relapsed Large Cell Carcinoma of the Lung
C0854977|T191|Relapsed Large Cell Carcinoma of Lung
CL446021|T061|Palliative Radiation Therapy for Metastatic Cancer
C1333986|T191|Hereditary Female Breast Carcinoma
C1333986|T191|Familial Female Breast Carcinoma
C0079380|T049|Frameshift Mutation
C0079380|T049|Out-of-Frame Mutations
C0079380|T049|Out of Frame Mutation
C0079380|T049|Frameshift Mutations
C0079380|T049|Frameshift Mutation function
C0079380|T049|Frameshift Mutation Abnormality
C0079380|T049|Mutations, Frameshift
C0079380|T049|frameshift mutation
C0079380|T049|Frame Shift Mutation
C0079380|T049|Out-of-Frame Mutation
C0079380|T049|frame-shift mutation
C0079380|T049|Mutation, Frame Shift
C0079380|T049|Mutations, Frame Shift
C0079380|T049|Frame Shift Mutations
C0079380|T049|Mutation, Out-of-Frame
C0079380|T049|Mutations, Out-of-Frame
C0079380|T049|Frameshift
C0079380|T049|Mutation, Frameshift
C0079380|T049|Reading Frame Shift Mutation
C0279644|T191|Childhood Acute Myelomonocytic Leukemia
C0279644|T191|myelomonoblastic leukemia, childhood acute
C0279644|T191|pediatric acute M4 leukemia
C0279644|T191|AMMoL, pediatric
C0279644|T191|Childhood Acute Myelomonocytic Leukemia (M4)
C0279644|T191|acute myelomonoblastic leukemia, childhood
C0279644|T191|M4 Pediatric Acute Myelomonocytic Leukemia
C0279644|T191|leukemia, childhood acute myelomonocytic
C0279644|T191|Pediatric AMMoL
C0279644|T191|childhood acute myelomonocytic leukemia
C0279644|T191|myelomonocytic leukemia, childhood acute
C0279644|T191|Pediatric AMML
C0279644|T191|AMML, pediatric
C0279644|T191|childhood AMML M4
C0279644|T191|Childhood AMMoL
C0279644|T191|Childhood Acute M4 Leukemia
C0279644|T191|M4 pediatric acute myelomonocytic leukemia
C0279644|T191|pediatric AMML
C0279644|T191|pediatric AMMoL
C0279644|T191|childhood acute M4 leukemia
C0279644|T191|M4 Childhood Acute Myelomonocytic Leukemia
C0279644|T191|M4 leukemia, childhood acute
C0279644|T191|AMMoL, childhood
C0279644|T191|AMML, childhood
C0279644|T191|childhood AMML
C0279644|T191|childhood acute myelomonocytic leukemia (M4)
C0279644|T191|pediatric acute myelomonocytic leukemia
C0279644|T191|Childhood AMML
C0279644|T191|Pediatric Acute Myelomonocytic Leukemia
C0279644|T191|acute myelomonocytic leukemia, childhood
C0279644|T191|Pediatric Acute M4 Leukemia
C0279644|T191|M4 childhood acute myelomonocytic leukemia
C0279644|T191|childhood AMMoL
C1706939|T061|Bilateral Prophylactic Oophorectomy
C0449454|T081|Stone size (observable entity)
C0449454|T081|Size of stone
C0449454|T081|Stone size
C1707605|T049|Cytosine to Guanosine Transversion Abnormality
C1707605|T049|Cytosine to Guanosine Transversion
C1707605|T049|Cytosine to Guanosine Mutation
C1300988|T201|Tumor size, largest metastasis, greatest dimension
C1300988|T201|Tumour size, largest metastasis, greatest dimension
C1300988|T201|Tumor size, largest metastasis, greatest dimension (observable entity)
C1332040|T191|AIDS-Related Cervical Carcinoma
C1332040|T191|AIDS-Related Uterine Cervix Carcinoma
C1332040|T191|AIDS-Related Cancer of Uterine Cervix
C1332040|T191|AIDS-related cervical cancer
C1332040|T191|AIDS-Related Cervical Cancer
C1332040|T191|AIDS Related Carcinoma of the Uterine Cervix
C1332040|T191|AIDS-Related Cancer of the Uterine Cervix
C1332040|T191|AIDS Related Carcinoma of Uterine Cervix
C1332040|T191|AIDS-Related Cervix Carcinoma
C1332040|T191|AIDS Related Cervical Cancer
C1332040|T191|AIDS-Related Uterine Cervix Cancer
C1334721|T033|Metastatic Mass
C0278846|T191|Invasive Malignant Thymoma
C0278846|T191|Thymoma Malignant Invasive
C0278846|T191|Thymoma malignant invasive
C0278846|T191|Malignant Thymoma, Invasive
C0862200|T191|Recurrent Mycosis Fungoides and Sezary Syndrome
C1333133|T191|Common Variant Anaplastic Large Cell Lymphoma
C1335938|T191|Secondary Chondrosarcoma
C2945767|T191|Childhood Malignant Liver Neoplasm
C2945767|T191|Pediatric Liver Cancer
C2945767|T191|Pediatric Cancer of Liver
C2945767|T191|Childhood Liver Cancer
C2945767|T191|liver cancer, childhood
C2945767|T191|Pediatric Cancer of the Liver
C2945767|T191|Liver cancer, child primary
C2945767|T191|childhood liver cancer
C2945767|T191|liver cancer, pediatric
C2945767|T191|pediatric liver cancer
C2945767|T191|Childhood Cancer of the Liver
C2945767|T191|Childhood Cancer of Liver
C0853968|T191|Recurrent Inflammatory Breast Carcinoma
C0853968|T191|Inflammatory carcinoma of breast recurrent
C0853968|T191|Recurrent Inflammatory Carcinoma of Breast
C0853968|T191|Recurrent Inflammatory Carcinoma of the Breast
C1512736|T191|Infiltrating Bladder Lymphoepithelioma-Like Carcinoma
C1384494|T191|Metastatic Carcinoma
C1384494|T191|Carcinoma, metastatic, NOS
C1384494|T191|Metastatic carcinoma
C1384494|T191|Secondary carcinoma
C1384494|T191|Carcinoma, metastatic
C1384494|T191|Carcinoma, metastatic (morphologic abnormality)
C1384494|T191|METASTATIC CARCINOMA
C0349656|T191|Spindle Cell (Sarcomatoid) Squamous Cell Skin Carcinoma
C0349656|T191|Spindle Cell Squamous Carcinoma of Skin
C0349656|T191|Spindle Cell Squamous Carcinoma of the Skin
C0279015|T061|Low-LET Implant Therapy
C0278810|T191|Localized Extrahepatic Bile Duct Carcinoma
C0278810|T191|bile duct cancer, localized extrahepatic
C0278810|T191|localized extrahepatic bile duct cancer
C0278810|T191|Localized Cancer of Extrahepatic Bile Duct
C0278810|T191|Localized Cancer of the Extrahepatic Bile Duct
C0278810|T191|Localized Extrahepatic Bile Duct Cancer
C0278810|T191|extrahepatic bile duct cancer, localized
C0684963|T191|Metastatic Malignant Neoplasm to the Pharynx
C0684963|T191|Metastatic Neoplasm to the Pharynx
C0684963|T191|Metastatic Tumor to the Pharynx
C0684963|T191|Metastasis to the Pharynx
C0220650|T191|Metastatic Malignant Neoplasm to the Brain
C0220650|T191|brain metastasis
C0220650|T191|Brain Metastasis
C0220650|T191|Metastases to brain parenchyma, NOS
C0220650|T191|Metast. to brain parenchyma, NOS
C0220650|T191|Metastatic Neoplasm to the Brain
C0220650|T191|Metastatic Tumor to the Brain
C0220650|T191|Brain Metastases
C1335520|T191|Acinar Prostate Adenocarcinoma, Signet Ring Variant
C1335520|T191|Signet Ring Cell Carcinoma of Prostate
C1335520|T191|Signet Ring Cell Carcinoma of the Prostate
C1335520|T191|Prostate Signet Ring Cell Carcinoma
C0684984|T191|Metastatic Malignant Neoplasm to the Larynx
C0684984|T191|Metastatic Tumor to the Larynx
C0684984|T191|Metastatic Neoplasm to the Larynx
C113813|T061|Involved Node Radiation Therapy
C113813|T061|INRT
C113813|T061|Involved node radiation therapy
C0334373|T191|Intraductal Papillary Adenocarcinoma with Invasion
C1334573|T191|Malignant Childhood Central Nervous System Neoplasm
C1334573|T191|Malignant Childhood Neoplasm of the Central Nervous System
C1334573|T191|Malignant Childhood Central Nervous System Neoplasms
C1334573|T191|Malignant Childhood Neoplasm of the CNS
C1334573|T191|Malignant Pediatric Central Nervous System Tumor
C1334573|T191|Childhood Malignant CNS Neoplasms
C1334573|T191|Malignant Pediatric CNS Neoplasm
C1334573|T191|Malignant Pediatric Tumor of CNS
C1334573|T191|Malignant Pediatric Tumor of Central Nervous System
C1334573|T191|Malignant Pediatric Central Nervous System Neoplasm
C1334573|T191|Malignant Central Nervous System Tumors of Childhood
C1334573|T191|Malignant Childhood Tumor of the CNS
C1334573|T191|Childhood Malignant Central Nervous System Tumors
C1334573|T191|Malignant Childhood Neoplasm of Central Nervous System
C1334573|T191|Childhood Malignant Central Nervous System Neoplasms
C1334573|T191|Malignant Childhood Tumor of CNS
C1334573|T191|Malignant Childhood Tumor of Central Nervous System
C1334573|T191|Malignant Pediatric Neoplasm of Central Nervous System
C1334573|T191|Childhood Malignant CNS Tumors
C1334573|T191|Malignant Pediatric Tumor of the Central Nervous System
C1334573|T191|Malignant Pediatric CNS Tumor
C1334573|T191|Malignant Central Nervous System Neoplasms of Childhood
C1334573|T191|Malignant Childhood CNS Neoplasm
C1334573|T191|Malignant Pediatric Neoplasm of the Central Nervous System
C1334573|T191|Malignant Childhood Central Nervous System Tumors
C1334573|T191|Malignant Childhood Tumor of the Central Nervous System
C1334573|T191|Malignant Pediatric Neoplasm of the CNS
C1334573|T191|Malignant Childhood Neoplasm of CNS
C1334573|T191|Malignant Pediatric Neoplasm of CNS
C1334573|T191|Malignant Pediatric Tumor of the CNS
C1334573|T191|Malignant Childhood Central Nervous System Tumor
C1334573|T191|Malignant Childhood CNS Tumor
C0238258|T191|Lymphangitic Carcinomatosis
C0238258|T191|Lymphangitis carcinomatosa (disorder)
C0238258|T191|LUNG, LYMPHANGITIC CANCER
C0238258|T191|LYMPHANGITIC CARCINOMATOSIS
C0238258|T191|Lymphangitis carcinomatosa
C0238258|T191|LYMPHANGITIS CARCINOMATOSIS
C0238258|T191|metastasis by lymphatic and interstitial infiltration
C0238258|T191|Lymphangitis carcinomatosis
C0238258|T191|LYMPHANGITIC METASTATIC DISEASE
C0238258|T191|lymphangitic carcinomatosis
C0854826|T191|Recurrent T-Cell Non-Hodgkin Lymphoma
C0854826|T191|Recurrent T-Cell and NK-Cell Non-Hodgkin's Lymphoma
C0854826|T191|T-Cell Lymphoma Relapsed
C0854826|T191|Recurrent T-Cell Lymphoma
C0854826|T191|Recurrent T-Cell Non-Hodgkin's Lymphoma
C0854826|T191|T-Cell Lymphoma Recurrent
C0854826|T191|Relapsed T-Cell Lymphoma
C2986562|T033|Spiculated Mass
C2986562|T033|stellate mass
C2986562|T033|irregular mass
C2986562|T033|spiculated mass
C2986562|T033|irregularly-shaped mass
C0280387|T191|Recurrent Nasopharyngeal Undifferentiated Carcinoma
C0280387|T191|Recurrent Nasopharyngeal Lymphoepithelioma
C0280387|T191|Nasopharyngeal lymphepithelioma recurrent
C0280387|T191|Relapsed Lymphoepithelioma of the Nasopharynx
C0280387|T191|Recurrent Lymphoepithelioma of Nasopharynx
C0280387|T191|nasopharyngeal lymphoepithelioma, recurrent
C0280387|T191|recurrent lymphoepithelioma of the nasopharynx
C0280387|T191|Relapsed Lymphoepithelioma of Nasopharynx
C0280387|T191|Relapsed Undifferentiated Carcinoma of Nasopharynx
C0280387|T191|Relapsed Nasopharyngeal Undifferentiated Carcinoma
C0280387|T191|Recurrent Lymphoepithelioma of the Nasopharynx
C0280387|T191|Relapsed Undifferentiated Carcinoma of the Nasopharynx
C0280387|T191|Nasopharyngeal lymphoepithelioma recurrent
C0280387|T191|Recurrent Undifferentiated Carcinoma of Nasopharynx
C0280387|T191|nasopharynx lymphoepithelioma, recurrent
C0280387|T191|Relapsed Nasopharyngeal Lymphoepithelioma
C0280387|T191|Recurrent Undifferentiated Carcinoma of the Nasopharynx
C0280387|T191|lymphoepithelioma of the nasopharynx, recurrent
C0549379|T191|Recurrent Malignant Neoplasm
C0549379|T191|Recurrent Malignant Tumor
C0549379|T191|recurrent cancer
C0549379|T191|Recurrent Cancer
C0549379|T191|Recurrent cancer
C0549379|T191|recurrence
C2919114|T034|Estrogen Receptor Status
C2919114|T034|ESTROGEN RECEPTOR STATUS
C2919114|T034|Estrogen receptor status (Z17)
C2919114|T034|Estrogen receptor status
C2919114|T034|ER Status
C2919114|T034|Encounter due to estrogen receptor status
C114836|T191|Recurrent Childhood Central Nervous System Embryonal Neoplasm
C1335718|T191|Recurrent Oral Cavity Carcinoma
C1335718|T191|Relapsed Oral Cavity Cancer
C1335718|T191|Recurrent Oral Cavity Cancer
C1335718|T191|Recurrent Carcinoma of the Oral Cavity
C1335718|T191|Recurrent Carcinoma of Mouth
C1335718|T191|Relapsed Mouth Carcinoma
C1335718|T191|Relapsed Carcinoma of Mouth
C1335718|T191|Recurrent Carcinoma of the Mouth
C1335718|T191|Recurrent Mouth Carcinoma
C1335718|T191|Relapsed Carcinoma of the Mouth
C1335718|T191|Relapsed Carcinoma of Oral Cavity
C1335718|T191|Relapsed Oral Cavity Carcinoma
C1335718|T191|Relapsed Carcinoma of the Oral Cavity
C1335718|T191|Recurrent Carcinoma of Oral Cavity
C0686031|T191|Metastatic Malignant Neoplasm to the Oropharynx
C0686031|T191|Metastasis to the Oropharynx
C0686031|T191|Metastatic Tumor to the Oropharynx
C0686031|T191|Metastatic Neoplasm to the Oropharynx
C481039|T116|Pertuzumab
C481039|T116|rhuMAb2C4
C481039|T116|Perjeta
C481039|T116|PERTUZUMAB
C481039|T116|rhuMAb 2C4
C481039|T116|pertuzumab
C481039|T116|2C4 Antibody
C481039|T116|monoclonal antibody 2C4
C481039|T116|2C4
C481039|T116|2C4 antibody
C481039|T116|MOAB 2C4
C481039|T116|Monoclonal Antibody 2C4
C481039|T116|rhuMAb-2C4
C481039|T116|MoAb 2C4
C1517577|T191|Invasive Mixed Breast Carcinoma
C1517577|T191|Infiltrating Mixed Breast Carcinoma
C1334184|T191|Infratentorial Glioblastoma
C1334184|T191|Infratentorial Glioblastoma Multiforme
C1334184|T191|Grade IV Infratentorial Astrocytic Tumor
C1334184|T191|Grade IV Infratentorial Astrocytic Neoplasm
C1332139|T191|Acinar Prostate Adenocarcinoma
C1332139|T191|Acinar Adenocarcinoma of Prostate
C1332139|T191|Prostatic Acinar Adenocarcinoma
C1332139|T191|Acinar Adenocarcinoma of the Prostate
C1519486|T191|Squamous Cell Breast Carcinoma, Large Cell Keratinizing Variant
C1333007|T191|Childhood Testicular Embryonal Carcinoma
C1333007|T191|Childhood Embryonal Carcinoma of the Testis
C1333007|T191|Pediatric Embryonal Carcinoma of the Testis
C1333007|T191|Childhood Embryonal Carcinoma of Testis
C1333007|T191|Pediatric Testicular Embryonal Carcinoma
C1333007|T191|Pediatric Embryonal Carcinoma of Testis
C2985552|T081|High-Dose-Rate Remote Brachytherapy
C2985552|T081|remote brachytherapy
C2985552|T081|high-dose-rate remote brachytherapy
C2985552|T081|high-dose-rate remote radiation therapy
C1705736|T116|Gene Fusion
C1705736|T116|fusion gene
C1705736|T116|Fusion gene in myxoid liposarcoma
C1705736|T116|Fusion, Gene
C1705736|T116|FUS/DDIT3 Fusion Protein
C1705736|T116|Fusions, Gene
C1705736|T116|FUS-CHOP protein fusion
C1705736|T116|TLS/CHOP Fusion Protein
C1705736|T116|FUS-DDIT3 Fusion Protein
C1705736|T116|RNA-Binding Protein FUS/DNA Damage-Inducible Transcript 3 Protein Fusion Protein
C1705736|T116|fus-like protein
C1705736|T116|TLS-CHOP Fusion Protein
C1705736|T116|fusion (involved in t(12;16) in malignant liposarcoma)
C1705736|T116|FUS-CHOP Fusion Protein
C1705736|T116|FUS
C1705736|T116|FUS/CHOP Fusion Protein
C1705736|T116|Gene Fusions
C1705736|T116|(AA).FUS.0
C1705736|T116|fusion, derived from t(12;16) malignant liposarcoma
C1705736|T116|Fusion Gene
C1705736|T116|fus/tls-chop oncogene
C1705736|T116|Gene Fusion Abnormality
C1333992|T191|Hereditary Ovarian Carcinoma
C1333992|T191|Familial Ovarian Carcinoma
C1300503|T201|Tumor size, dominant nodule, greatest dimension, in specimen obtained by radical prostatectomy
C1300503|T201|Tumour size, dominant nodule, greatest dimension, in specimen obtained by radical prostatectomy
C1300503|T201|Tumor size, dominant nodule, greatest dimension, in specimen obtained by radical prostatectomy (observable entity)
C1332056|T191|AIDS-Related Plasmablastic Lymphoma of Mucosa Site
C0162505|T061|Boron Neutron Capture Therapy
C0162505|T061|boron neutron capture therapy
C0162505|T061|THER BORON NEUTRON CAPTURE
C0162505|T061|Therapy, Boron Neutron Capture
C0162505|T061|Neutron Capture Therapy, Boron
C0162505|T061|Therapy, Boron-Neutron Capture
C0162505|T061|NEUTRON CAPTURE THER BORON
C0162505|T061|Boron-Neutron Capture Therapy
C0162505|T061|BNCT
C0162505|T061|BORON NEUTRON CAPTURE THER
C0851238|T061|Lumpectomy
C0851238|T061|Lumpectomy of breast
C0851238|T061|Breast lump removal
C0851238|T061|Limited Resection Mastectomies
C0851238|T061|Limited Resection Mastectomy
C0851238|T061|Mastectomy, Local Excision
C0851238|T061|Local Excision Mastectomy
C0851238|T061|Tylectomy of breast
C0851238|T061|Mastectomies, Limited Resection
C0851238|T061|Breast lump removal NOS
C0851238|T061|Resection Mastectomy, Limited
C0851238|T061|Partial Mastectomy
C0851238|T061|Lumpectomy of Breast
C0851238|T061|Excision Mastectomies, Local
C0851238|T061|Lumpectomy of breast (procedure)
C0851238|T061|Mastectomies, Local Excision
C0851238|T061|Tylectomy (procedure)
C0851238|T061|Resection Mastectomies, Limited
C0851238|T061|partial mastectomy
C0851238|T061|Excision of breast lump
C0851238|T061|Breast lumpectomy
C0851238|T061|Tylectomy
C0851238|T061|lumpectomy
C0851238|T061|Mastectomy, Limited Resection
C0851238|T061|Excision Mastectomy, Local
C0851238|T061|Local Excision Mastectomies
C1327920|T191|Childhood Chronic Myelogenous Leukemia, BCR-ABL1 Positive
C1327920|T191|Childhood Chronic Myelogenous Leukemia
C1327920|T191|Childhood Chronic Myeloid Leukemia
C1327920|T191|Childhood CML
C0279636|T191|Childhood Acute Myeloid Leukemia with Maturation
C0279636|T191|Childhood Acute Myeloblastic Leukemia with Maturation (M2)
C0279636|T191|M2 Pediatric Acute Granulocytic Leukemia with Maturation
C0279636|T191|M2 Pediatric Acute Myeloid Leukemia with Maturation
C0279636|T191|Childhood Acute Granulocytic Leukemia with Maturation
C0279636|T191|M2 Childhood Acute Myelogenous Leukemia with Maturation
C0279636|T191|Pediatric Acute Myeloblastic Leukemia with Maturation
C0279636|T191|Pediatric Acute Granulocytic Leukemia with Maturation
C0279636|T191|Pediatric Acute Myelocytic Leukemia with Maturation
C0279636|T191|Pediatric Acute M2 Leukemia
C0279636|T191|M2 Pediatric Acute Myeloblastic Leukemia with Maturation
C0279636|T191|Childhood Acute Myelocytic Leukemia with Maturation
C0279636|T191|M2 Pediatric AGL
C0279636|T191|M2 Pediatric Acute Myelogenous Leukemia
C0279636|T191|Childhood Acute Myeloblastic Leukemia with Maturation
C0279636|T191|Pediatric AGL with Maturation
C0279636|T191|M2 Childhood Acute Myelocytic Leukemia with Maturation
C0279636|T191|M2 Childhood Acute Myelogenous Leukemia
C0279636|T191|Childhood Acute Myelogenous Leukemia with Maturation
C0279636|T191|M2 Pediatric Acute Myelocytic Leukemia with Maturation
C0279636|T191|Pediatric Acute Myeloid Leukemia with Maturation
C0279636|T191|Childhood Acute M2 Leukemia
C0279636|T191|M2 Childhood Acute Myeloblastic Leukemia with Maturation
C0279636|T191|M2 Childhood AGL
C0279636|T191|M2 Pediatric Acute Myelogenous Leukemia with Maturation
C0279636|T191|Pediatric Acute Myelogenous Leukemia with Maturation
C0279636|T191|M2 Childhood Acute Myeloid Leukemia with Maturation
C1708262|T049|Guanosine to Cytosine Transversion Abnormality
C1708262|T049|Guanosine to Cytosine Transversion
C1708262|T049|Guanosine to Cytosine Mutation
C1335425|T191|Plasma Cell Myeloma Post-Transplant Lymphoproliferative Disorder
C1335425|T191|Plasma Cell Myeloma PTLD
C0279759|T034|Progesterone Receptor Positive
C0279759|T034|PR+
C0279759|T034|positive progesterone receptor
C0279759|T034|progesterone receptor positive
C0221783|T033|Vaginal Mass
C0221783|T033|VAGINAL MASS
C0221783|T033|Vaginal mass (finding)
C0221783|T033|Vaginal mass
C0238869|T033|Buttock Mass
C0238869|T033|BUTTOCK MASS
C1334463|T191|Lymphohistiocytic Variant Anaplastic Large Cell Lymphoma
CL414408|T191|Childhood Glioblastoma
CL414408|T191|Brain tumor, child: Glioblastoma
CL414408|T191|grade IV childhood astrocytic neoplasm
CL414408|T191|Grade IV Childhood Astrocytic Tumor
CL414408|T191|Grade IV Pediatric Astrocytic Neoplasm
CL414408|T191|pediatric glioblastoma multiforme
CL414408|T191|glioblastoma multiforme, childhood
CL414408|T191|Grade IV Childhood Astrocytic Neoplasm
CL414408|T191|Pediatric Glioblastoma Multiforme
CL414408|T191|grade IV childhood astrocytic tumor
CL414408|T191|Grade IV Pediatric Astrocytic Tumor
CL414408|T191|grade IV childhood astrocytoma
CL414408|T191|grade IV pediatric astrocytic tumor
CL414408|T191|Childhood Glioblastoma Multiforme
CL414408|T191|grade IV pediatric astrocytic neoplasm
CL414408|T191|astrocytoma, grade IV childhood
CL414408|T191|childhood glioblastoma
CL414408|T191|childhood glioblastoma multiforme
C1332987|T191|Childhood Ovarian Choriocarcinoma
C1332987|T191|Pediatric Choriocarcinoma of the Ovary
C1332987|T191|Childhood Choriocarcinoma of the Ovary
C1332987|T191|Pediatric Ovarian Choriocarcinoma
C1332987|T191|Pediatric Choriocarcinoma of Ovary
C1332987|T191|Childhood Choriocarcinoma of Ovary
C0677861|T191|Bilateral Malignant Neoplasm
C0677861|T191|Bilateral Cancer
C0677861|T191|Bilateral Malignant Tumor
C0948840|T191|Meningeal Leukemia
C0948840|T191|Meningeal leukemia
C0948840|T191|meningitis, leukemic
C0948840|T191|meningeal leukemia
C0948840|T191|leptomeningitis, leukemic
C0948840|T191|leukemic meningitis
C0948840|T191|Meningeal leukaemia
C0948840|T191|Leukemic Leptomeningitis
C0948840|T191|Leukemic Meningitis
C0948840|T191|leukemic leptomeningitis
C0677726|T191|Recurrent Aggressive Adult Non-Hodgkin Lymphoma
C0677726|T191|Aggressive Recurrent Adult Non-Hodgkin's Lymphoma
C0677726|T191|Recurrent Aggressive Adult Non-Hodgkin's Lymphoma
C0677726|T191|Recurrent Adult Aggressive Non-Hodgkin's Lymphoma
C1332550|T033|Bilateral Mass
C0686377|T191|Metastatic Malignant Neoplasm to the Central Nervous System
C0686377|T191|CNS Metastasis
C0686377|T191|Metastatic Neoplasm to the Central Nervous System
C0686377|T191|Metastatic Tumor to the CNS
C0686377|T191|Central Nervous System Metastasis
C0686377|T191|central nervous system metastasis
C0686377|T191|Metastatic Neoplasm to the CNS
C0686377|T191|Metastatic Tumor to the Central Nervous System
C0686377|T191|Central Nervous System Metastases
C0686377|T191|CNS Metastases
C0686377|T191|CNS metastasis
C0279567|T191|Paget Disease of the Breast with Invasive Ductal Carcinoma
C0279567|T191|Paget's Disease and Invasive Ductal Carcinoma of the Breast
C0279567|T191|Paget's Disease and Infiltrating Ductal Carcinoma of Breast
C0279567|T191|Paget's Disease of Breast with Infiltrating Ductal Carcinoma
C0279567|T191|Paget's Disease of the Breast with Invasive Ductal Carcinoma
C0279567|T191|Paget's Disease of the Breast with Infiltrating Ductal Carcinoma
C0279567|T191|Paget's Disease and Invasive Ductal Carcinoma of Breast
C0279567|T191|Paget's Disease of Breast with Invasive Ductal Carcinoma
C0279567|T191|Paget's Disease and Infiltrating Ductal Carcinoma of the Breast
C1332941|T191|Childhood Acute Monoblastic and Monocytic Leukemia
C1332941|T191|Childhood Acute Monoblastic Leukemia and Acute Monocytic Leukemia
C1332941|T191|Childhood Acute Monoblastic and Monocytic Leukemia (M5)
C1512737|T191|Infiltrating Bladder Urothelial Carcinoma, Clear Cell Variant
C0547070|T061|Ablation Therapy
C0547070|T061|Ablation
C0547070|T061|ablation
C0547070|T061|ablate
C0547070|T061|ABLATION
C0547070|T061|ablat
C0547070|T061|Ablation - action (qualifier value)
C0547070|T061|Ablation - action
C1516197|T049|Cancer Gene Mutation
C1883578|T121|Xinidamine
C1883578|T121|XINIDAMINE
C1883578|T121|1-(2,4-Dimethylbenzyl)-1H-indazole-3-carboxylic Acid
C113811|T061|Extended-Field Radiation Therapy
C113811|T061|Extended field radiation
C113811|T061|EFRT
C1300495|T201|Tumor size, dominant nodule, additional dimension
C1300495|T201|Tumor size, dominant nodule, additional dimension (observable entity)
C1300495|T201|Tumour size, dominant nodule, additional dimension
C1332955|T191|Childhood Central Nervous System Mature Teratoma
C1300498|T201|Tumor size, dominant nodule, in specimen obtained by prostatic enucleation
C1300498|T201|Tumour size, dominant nodule, in specimen obtained by prostatic enucleation
C1300498|T201|Tumor size, dominant nodule, in specimen obtained by prostatic enucleation (observable entity)
C0475392|T185|Tumor stage T3bi
C0475392|T185|Tumour stage T3bi
C0475392|T185|Tumor stage T3bi (finding)
C2985439|T049|de novo Mutation
C2985439|T049|de novo mutation
C2985439|T049|new mutation
C1883035|T033|Single Cell Necrosis
C1337019|T191|Well Differentiated Malignant Neoplasm
C1332996|T191|Childhood B Lymphoblastic Lymphoma
C1332996|T191|Childhood B-Lymphoblastic Lymphoma
C1332996|T191|Childhood Precursor B-Lymphoblastic Lymphoma
C0424863|T033|Length of lump
C0424863|T033|Length of lump (observable entity)
C1517030|T061|Extensive Radiation
C0278773|T191|Localized Non-Resectable Adult Liver Carcinoma
C0278773|T191|Localized Unresectable Adult Primary Cancer of Liver
C0278773|T191|Localized Unresectable Adult Primary Cancer of the Liver
C0278773|T191|Localized Unresectable Adult Liver Carcinoma
C0278773|T191|Localized Unresectable Adult Primary Liver Cancer
C0278773|T191|Localized Non-Resectable Adult Liver Cancer
C1332957|T191|Childhood Central Nervous System Primitive Neuroectodermal Tumor
C1332957|T191|Childhood CNS Primitive Neuroectodermal Tumor
C1332957|T191|Pediatric CNS PNET
C1332957|T191|Childhood CNS PNET
C1332957|T191|Pediatric CNS Primitive Neuroectodermal Neoplasm
C1332957|T191|Pediatric Central Nervous System Primitive Neuroectodermal Neoplasm
C1332957|T191|Pediatric Central Primitive Neuroectodermal Neoplasm
C1332957|T191|Childhood CNS Primitive Neuroectodermal Neoplasm
C1332957|T191|Pediatric Central Primitive Neuroectodermal Tumor
C1332957|T191|Childhood Central Primitive Neuroectodermal Neoplasm
C1332957|T191|Childhood Central Primitive Neuroectodermal Tumor
C1332957|T191|Childhood Central Nervous System PNET
C1332957|T191|Pediatric CNS Primitive Neuroectodermal Tumor
C1332957|T191|Pediatric Central Nervous System Primitive Neuroectodermal Tumor
C1332957|T191|Childhood Central Nervous System Primitive Neuroectodermal Neoplasm
C0445080|T033|N2b Stage Finding
C0445080|T033|N2b Lymph Node Finding
C0445080|T033|N2b Node Finding
C0445080|T033|N2b Lymph Node Stage
C0445080|T033|N2b Node Stage
C0445080|T033|Lymph Node Stage N2b
C0445080|T033|N2b Stage
C0445080|T033|N2b Cancer Stage Finding
C0445080|T033|N2b
C0445080|T033|Node Stage N2b
C0445080|T033|Node stage N2b
C0445080|T033|N2b TNM Finding
C0445080|T033|N2b Regional Lymph Node Stage Finding
C0445080|T033|N2b Regional Lymph Nodes Finding
C0445080|T033|Node stage N2b (finding)
C0431108|T191|Anaplastic Oligoastrocytoma
C0431108|T191|Anaplastic oligoastrocytoma
C0431108|T191|Anaplastic Mixed Glioma
C0431108|T191|anaplastic oligoastrocytoma (WHO grade III)
C0431108|T191|WHO Grade III Mixed Glioma
C0431108|T191|anaplastic oligoastrocytoma
C0431108|T191|Anaplastic oligoastrocytoma (morphologic abnormality)
C0279984|T191|Childhood Liposarcoma
C0279984|T191|pediatric liposarcoma
C0279984|T191|liposarcoma, pediatric
C0279984|T191|childhood liposarcoma
C0279984|T191|liposarcoma, childhood
C0279984|T191|Pediatric Liposarcoma
C0279984|T191|sarcoma, lipo-, childhood
C0347015|T191|Metastatic Malignant Neoplasm to the Pituitary Gland
C0347015|T191|Metastatic Neoplasm to the Pituitary Gland
C0347015|T191|Metastasis to Pituitary Gland
C1302530|T191|Prostate Squamous Cell Carcinoma
C1302530|T191|Squamous cell carcinoma of prostate (disorder)
C1302530|T191|Squamous Cell Carcinoma of Prostate
C1302530|T191|Squamous Cell Carcinoma of the Prostate
C1302530|T191|Squamous cell carcinoma of prostate
C1512750|T191|Infiltrating Renal Pelvis and Ureter Urothelial Carcinoma
C1512750|T191|Infiltrating Renal Pelvis and Ureter Transitional Cell Carcinoma
C0457422|T033|V1 stage
C0457422|T033|Venous Stage V1
C0457422|T033|V1 TNM Finding
C0457422|T033|V1 Stage Finding
C0457422|T033|V1
C0457422|T033|V1 stage (finding)
C0457422|T033|V1: microscopic venous invasion
C0457422|T033|V1 Venous Invasion Finding
C0457422|T033|V1 Stage
C0457422|T033|V1 Cancer Stage Finding
C0457422|T033|Venous stage V1
C0457422|T033|V1 Venous Stage
C0475396|T185|T4b Stage Finding
C0475396|T185|Tumour stage T4b
C0475396|T185|Tumor stage T4b
C0475396|T185|T4b Primary Tumor Stage Finding
C0475396|T185|T4b Primary Tumor Finding
C0475396|T185|T4b Stage
C0475396|T185|T4b TNM Finding
C0475396|T185|Tumor stage T4b (finding)
C0475396|T185|T4b tumor stage
C0475396|T185|T4b
C0475396|T185|T4b Tumor Finding
C0475396|T185|T4b Tumor Stage
C0475396|T185|T4b Cancer Stage Finding
C0475396|T185|Tumor Stage T4b
C0014859|T191|Esophageal Mass
C0014859|T191|Esophageal tumor
C0014859|T191|Esophageal neoplasm NOS
C0014859|T191|Neoplasm of esophagus
C0014859|T191|Esophagus Neoplasms
C0014859|T191|Esophageal mass
C0014859|T191|Oesophageal neoplasm
C0014859|T191|Neoplasm of oesophagus
C0014859|T191|esophagus neoplasm
C0014859|T191|Neoplasm of Esophagus
C0014859|T191|Tumor of the Esophagus
C0014859|T191|ESOPHAGUS NEOPL
C0014859|T191|Esophageal Neoplasm
C0014859|T191|Esophageal Neoplasms
C0014859|T191|Oesophageal neoplasm NOS
C0014859|T191|esophageal neoplasm
C0014859|T191|Tumor of Esophagus
C0014859|T191|Neoplasm, Esophagus
C0014859|T191|Oesophageal mass
C0014859|T191|Tumor of esophagus
C0014859|T191|esophageal tumor or cancer
C0014859|T191|ESOPHAGEAL TUMOR
C0014859|T191|Esophagus Tumor
C0014859|T191|Neoplasms, Esophagus
C0014859|T191|Neoplasm, Esophageal
C0014859|T191|NEOPL ESOPHAGEAL
C0014859|T191|Tumour of oesophagus
C0014859|T191|Esophageal mass (finding)
C0014859|T191|Neoplasm of the Esophagus
C0014859|T191|Esophageal Neoplasms, Benign and Malignant
C0014859|T191|Oesophageal Mass
C0014859|T191|Esophageal Tumor
C0014859|T191|Esophageal neoplasm
C0014859|T191|Neoplasms, Esophageal
C0014859|T191|ESOPHAGEAL NEOPL
C0014859|T191|Esophageal Neoplasms [Disease/Finding]
C0014859|T191|Neoplasm of esophagus (disorder)
C0014859|T191|Esophageal Tumors
C0014859|T191|esophageal cancer
C0014859|T191|Esophagus Neoplasm
C0279650|T191|Childhood Acute Megakaryoblastic Leukemia
C0279650|T191|Pediatric Acute Megakaryocytic Leukemia
C0279650|T191|Pediatric Acute M7 Leukemia
C0279650|T191|Childhood Acute M7 Leukemia
C0279650|T191|leukemia, childhood acute megakaryocytic
C0279650|T191|M7 Childhood Acute Megakaryocytic Leukemia
C0279650|T191|Childhood Acute Megakaryocytic Leukemia
C0279650|T191|Pediatric Acute Megakaryoblastic Leukemia
C0279650|T191|M7 Pediatric Acute Megakaryocytic Leukemia
C0279650|T191|pediatric acute megakaryocytic leukemia
C0279650|T191|childhood acute megakaryocytic leukemia (M7)
C0279650|T191|megakaryocytic leukemia, childhood acute
C0279650|T191|acute megakaryocytic leukemia, childhood
C0279650|T191|M7 pediatric acute megakaryocytic leukemia
C0279650|T191|M7 childhood acute megakaryocytic leukemia
C0279650|T191|Childhood Acute Megakaryocytic Leukemia (M7)
C1335458|T191|Postsurgical Stage III Hepatoblastoma
C1882498|T061|Proton Beam Radiation Therapy
C1882498|T061|proton beam radiation therapy
C1336860|T191|Undifferentiated Malignant Neoplasm
C0279914|T191|Stage II Childhood Hodgkin Lymphoma
C0279914|T191|Pediatric Hodgkin's Lymphoma Stage II
C0279914|T191|Stage II Pediatric Hodgkin's Lymphoma
C0279914|T191|Childhood Hodgkin's Lymphoma Stage II
C0279914|T191|Pediatric Hodgkin's Disease Stage II
C0279914|T191|Stage II Childhood Hodgkin's Lymphoma
C0279914|T191|Childhood Hodgkin's Disease Stage II
C0279914|T191|stage II childhood Hodgkin lymphoma
C1299212|T201|Polyp size
C1299212|T201|Polyp size (observable entity)
C0475276|T081|Tumor Volume
C0475276|T081|Tumor volume (observable entity)
C0475276|T081|Tumour volume
C0475276|T081|Tumor volume
C0475276|T081|tumor volume
C0475276|T081|Volume, Tumor
C0347014|T191|Metastatic Malignant Neoplasm to the Nervous System
C0347014|T191|Metastasis to the Nervous System
C0347014|T191|Secondary Malignant Neoplasm to the Nervous System
C0347014|T191|Metastatic Neoplasm to the Nervous System
C0347014|T191|Secondary Malignant Tumor to the Nervous System
C0347014|T191|Metastatic Tumor to the Nervous System
C0347014|T191|Metastases to Nervous System
C1511304|T191|Breast Carcinoma with Osteoclastic Giant Cells
C1335491|T191|Primary Systemic Anaplastic Large Cell Lymphoma, ALK-Negative
C1335491|T191|Primary Systemic ALK-Negative Anaplastic Large Cell Lymphoma
C1515107|T191|Synchronous Bilateral Breast Carcinoma
C2983137|T191|Colon Carcinoma Metastatic to the Lung
C1879499|T061|AC-T-T Regimen
C1879499|T061|AC-T-T regimen
C1879499|T061|AC-T-T
C1879499|T061|AC-TH regimen
C1879499|T061|sequential AC/Taxol-Trastuzumab regimen
C1879499|T061|Sequential AC/Taxol-Trastuzumab Regimen
C0334233|T191|Pleomorphic Carcinoma
C0334233|T191|Pleomorphic carcinoma
C0334233|T191|Pleomorphic carcinoma (morphologic abnormality)
C1377767|T191|Recurrent Malignant Nasopharyngeal Neoplasm
C1377767|T191|Malignant neoplasm of nasopharynx recurrent
C1377767|T191|Malignant nasopharyngeal neoplasm recurrent
C0855085|T191|Recurrent Nodular Sclerosis Classical Hodgkin Lymphoma
C0855085|T191|Recurrent Hodgkin's Nodular Sclerosis
C0855085|T191|Recurrent Nodular Sclerosis Hodgkin's Lymphoma
C0855085|T191|Relapsed Nodular Sclerosis Hodgkin's Disease
C0855085|T191|Hodgkin's disease nodular sclerosis recurrent
C0855085|T191|Relapsed Nodular Sclerosis Hodgkin's Lymphoma
C0855085|T191|Recurrent Nodular Sclerosis Hodgkin's Disease
C0855085|T191|Recurrent Nodular Sclerosis Hodgkin Lymphoma
C1512413|T034|Her2/Neu Status
C1512413|T034|ERBB2 Status
C1512413|T034|Her2/Neu Value
C1332042|T191|AIDS-Related Diffuse Large B-cell Lymphoma
C3275043|T061|Ablation of Cardiac Accessory Pathway
C3275043|T061|ABLATION, ACCESSORY PATHWAYS
C1517579|T191|Infiltrating Bladder Urothelial Carcinoma, Micropapillary Variant
C0449457|T082|Nodule size
C0449457|T082|Nodule size (observable entity)
C0449457|T082|Size of nodule
C0746921|T047|Lymph Node Mass
C0746921|T047|Nodal Mass
C1512743|T191|Infiltrating Bladder Urothelial Carcinoma Sarcomatoid Variant
C116429|T061|3-Dimensional Ultrasound-Guided Radiation Therapy
C116429|T061|3D Ultrasound-Guided Radiation Therapy
C1334006|T191|High Grade Mucoepidermoid Breast Carcinoma
C1334006|T191|High-Grade Mucoepidermoid Carcinoma of the Breast
C1334006|T191|High-Grade Mucoepidermoid Carcinoma of Breast
C1334543|T191|Macrotrabecular Hepatoblastoma
C1711391|T191|Recurrent Adult Hepatocellular Carcinoma
C0346993|T191|Metastatic Malignant Neoplasm to the Breast
C0346993|T191|Metastatic Neoplasm to the Breast
C0346993|T191|Metastatic Tumor to the Breast
C0346993|T191|Metastatic Cancer to the Breast
C0346993|T191|Breast Metastasis
C0346993|T191|Breast Metastases
CL448471|T191|Metastatic Carcinoma to the Lung
C1514496|T061|Prophylactic Cranial Irradiation
C1514496|T061|PCI
C1514496|T061|prophylactic cranial irradiation
C1882994|T061|Selective External Radiation Therapy
C1882994|T061|SERT
C1882994|T061|selective external radiation therapy
C0246415|T121|Docetaxel
C0246415|T121|[2aR-[2a alphaa,4beta,4a beta,6beta,9alpha,(alphaR*,betaS*),-11alpha,12alpha,12a alpha,12b alpha]]-beta-[[(1,1-dimethylethoxy)carbonyl]-amino]-alpha-hydroxybenzemepropanoic Acid 12b-(Acetyloxy)-12(benzyloxy)-2a,3,4,4a,5,6,8,10,11,12,12a,12b-dodecahydeo-4,-6,11-trihydroxy-4a,8,13,13-tetramethyl-5-oxo-7,11-methano-1H-cyclodeca[3,4]benz[1,2-b]oxet-9-yl Ester
C0246415|T121|N-Debenzoyl-N-(tert-butoxycarbonyl)-10-deacetyltaxol
C0246415|T121|Taxotere
C0246415|T121|[2aR-[2a alphaa,4beta,4a beta,6beta,9alpha,(alphaR*,betaS*),-11alpha,12alpha,12a alpha,12b alpha]]-beta-[[(1,1-dimethylethoxy)carbonyl]-amino]-alpha-hydroxybenzemepropanoic acid 12b-(Acetyloxy)-12(benzyloxy)-2a,3,4,4a,5,6,8,10,11,12,12a,12b-dodecahydeo-4,-6,11-trihydroxy-4a,8,13,13-tetramethyl-5-oxo-7,11-methano-1H-cyclodeca[3,4]benz[1,2-b]oxet-9-yl ester
C0246415|T121|Docetaxel (product)
C0246415|T121|628503
C0246415|T121|RP 56976
C0246415|T121|RP56976
C0246415|T121|Benzenepropanoic acid, beta-(((1,1-dimethylethoxy)carbonyl)amino)-alpha-hydroxy-, 12b-(acetyloxy)-12-(benzoyloxy)-2a,3,4,4a,5,6,9,10,11,12,12a,12b-dodecahydro-4,6,11-trihydroxy-4a,8,13,13-tetramethyl-5-oxo-7,11-methano-1H-cyclodeca(3,4)benz(1,2-b)oxet-9-y
C0246415|T121|docetaxol
C0246415|T121|docetaxel
C0246415|T121|Benzenepropanoic acid, beta-(((1,1-dimethylethoxy)carbonyl)amino)-alpha-hydroxy-, 12b-(acetyloxy)-12-(benzoyloxy)-2a,3,4,4a,5,6,9,10,11,12,12a,12b-dodecahydro-4,6,11-trihydroxy-4a,8,13,13-tetramethyl-5-oxo-7,11-methano-1H-cyclodeca(3,4)benz(1,2-b)oxet-9-yl ester
C0246415|T121|40466
C0246415|T121|Taxotere Injection Concentrate
C0246415|T121|taxotere
C0246415|T121|DOCEtaxel
C0246415|T121|TXT
C0246415|T121|DOCETAXEL
C0246415|T121|N-debenzoyl-N-(tert-butoxycarbonyl)-10-deacetyltaxol
C0246415|T121|114977-28-5
C0246415|T121|Docetaxel (substance)
C0246415|T121|docetaxel [Chemical/Ingredient]
C0246415|T121|N-debenzoyl-N-tert-butoxycarbonyl-10-deacetyltaxol
C1512749|T191|Infiltrating Bladder Urothelial Carcinoma with Trophoblastic Differentiation
C0279999|T191|Recurrent Adult Non-Hodgkin Lymphoma
C0279999|T191|Adult Recurrent Non-Hodgkin's Lymphoma
C0279999|T191|Relapsed Adult Non-Hodgkin's Lymphoma
C0279999|T191|Recurrent Adult Non-Hodgkin's Lymphoma
C0279999|T191|Adult Relapsed Non-Hodgkin's Lymphoma
CL448459|T191|Recurrent Malignant Hypopharyngeal Neoplasm
C2348970|T061|High-Intensity Focused Ultrasound Ablation
C2348970|T061|HIFU
C2348970|T061|high-intensity focused ultrasound therapy
C1367872|T191|Metastatic Neoplasm of the Ureter
C1367872|T191|Metastatic Neoplasm of Ureter
C1367872|T191|Ureter Metastatic Malignant Neoplasm
C0279018|T061|High-LET Pion Therapy
C0279018|T061|therapy, high-LET pion
C0334590|T191|Anaplastic Oligodendroglioma
C0334590|T191|Oligodendrogliomas, Anaplastic
C0334590|T191|WHO Grade III Oligodendroglial Tumor
C0334590|T191|UNDIFFERENTIATED OLIGODENDROGLIOMA
C0334590|T191|anaplastic oligodendroglioma (WHO grade III)
C0334590|T191|WHO GRADE III OLIGODENDROGLIAL TUMOR
C0334590|T191|MALIGNANT OLIGODENDROGLIOMA
C0334590|T191|Anaplastic oligodendroglioma
C0334590|T191|Oligodendroglioma, anaplastic
C0334590|T191|Anaplastic Oligodendrogliomas
C0334590|T191|Oligodendroglioma, Malignant
C0334590|T191|Oligodendroglioma, Anaplastic
C0334590|T191|Oligodendroglioma malignant
C0334590|T191|OLIGODENDROGLIOMA
C0334590|T191|anaplastic oligodendroglioma
C0334590|T191|Oligodendroglioma, anaplastic (morphologic abnormality)
C0334590|T191|Malignant oligodendroglioma
C0334590|T191|WHO Grade III Oligodendroglial Neoplasm
C0334590|T191|OLIGODENDROGLIOMA, ANAPLASTIC, MALIGNANT
C0334590|T191|MALIGNANT
C0334590|T191|WHO GRADE III OLIGODENDROGLIAL NEOPLASM
C0334590|T191|Undifferentiated Oligodendroglioma
C0334590|T191|Malignant Oligodendroglioma
C1831994|T061|Selective Internal Radiation Therapy
C1831994|T061|SIRT
C1831994|T061|selective internal radiation therapy
C1332281|T191|Anaplastic Diencephalic Astrocytoma
C1332281|T191|Grade III Diencephalic Astrocytic Neoplasm
C1332281|T191|Grade III Astrocytoma of Diencephalon
C1332281|T191|Undifferentiated Astrocytoma of the Diencephalon
C1332281|T191|Undifferentiated Astrocytoma of Diencephalon
C1332281|T191|Diencephalic Anaplastic Astrocytoma
C1332281|T191|Anaplastic Astrocytoma of the Diencephalon
C1332281|T191|Grade III Astrocytic Neoplasm of the Diencephalon
C1332281|T191|Grade III Astrocytic Neoplasm of Diencephalon
C1332281|T191|Grade III Diencephalic Astrocytoma
C1332281|T191|Grade III Diencephalic Astrocytic Tumor
C1332281|T191|Anaplastic Astrocytoma of Diencephalon
C1332281|T191|Undifferentiated Diencephalic Astrocytoma
C1332281|T191|Grade III Astrocytic Tumor of Diencephalon
C1332281|T191|Grade III Astrocytic Tumor of the Diencephalon
C1332281|T191|Grade III Astrocytoma of the Diencephalon
C1300501|T201|Tumor size, dominant nodule, additional dimension, in specimen obtained by radical prostatectomy
C1300501|T201|Tumor size, dominant nodule, additional dimension, in specimen obtained by radical prostatectomy (observable entity)
C1300501|T201|Tumour size, dominant nodule, additional dimension, in specimen obtained by radical prostatectomy
C1335702|T191|Recurrent Gastrointestinal Carcinoma
C1335702|T191|Recurrent Gastrointestinal System Carcinoma
C1335702|T191|Recurrent Gastrointestinal System Cancer
C1711210|T033|Cancer stage
C1711210|T033|Generic TNM Finding
C1708231|T033|Generic Primary Tumor TNM Finding
C1334747|T191|Methotrexate-Associated Follicular Lymphoma
C0862489|T191|Metastatic Endometrial Adenocarcinoma
C0862489|T191|Endometrial adenocarcinoma metastatic
C0862489|T191|Adenocarcinoma endometrial metastatic
C1706718|T049|Adenosine to Thymidine Transversion Abnormality
C1706718|T049|Adenosine to Thymidine Mutation
C1706718|T049|Adenosine to Thymidine Transversion
C0334496|T191|Intracanalicular Fibroadenoma
C0334496|T191|Intracanalicular Fibroadenoma of the Breast
C0334496|T191|Intracanalicular Fibroadenoma of Breast
C0334496|T191|Intracanalicular fibroadenoma
C0334496|T191|Intracanalicular Breast Fibroadenoma
C0334496|T191|BREAST, FIBROADENOMA, INTRACANALICULAR
C0334496|T191|Intracanalicular fibroadenoma (morphologic abnormality)
C0279565|T191|Invasive Lobular Breast Carcinoma
C0279565|T191|Invasive Lobular Carcinoma
C0279565|T191|Infiltrating Lobular Breast Carcinoma
C0279565|T191|invasive lobular breast carcinoma
C0279565|T191|lobular invasive breast carcinoma
C0279565|T191|Infiltrating lobular carcinoma, NOS
C0279565|T191|Invasive Lobular Carcinoma of the Breast
C0279565|T191|Infiltrating Lobular Adenocarcinoma
C0279565|T191|Invasive Lobular Carcinoma of Breast
C0279565|T191|Invasive lobular breast carcinoma
C0279565|T191|Invasive Lobular Carcinoma, Classic Type
C0279565|T191|Lobular breast carcinoma invasive
C0279565|T191|Classic Invasive Lobular Carcinoma
C0279565|T191|Infiltrating Lobular Carcinoma of Breast
C0279565|T191|Invasive Lobular Adenocarcinoma
C0279565|T191|Infiltrating Lobular Carcinoma of the Breast
C0281708|T191|Recurrent Childhood Burkitt Lymphoma
C0281708|T191|recurrent small noncleaved cell lymphoma, childhood
C0281708|T191|relapsed childhood small noncleaved cell lymphoma
C0281708|T191|pediatric small noncleaved cell lymphoma, relapsed
C0281708|T191|recurrent childhood small noncleaved cell lymphoma
C0281708|T191|small noncleaved cell lymphoma, childhood, relapsed
C0281708|T191|lymphoma, recurrent childhood small noncleaved cell
C0281708|T191|Recurrent Childhood Small Non-Cleaved Cell Lymphoma
C0281708|T191|lymphoma, relapsed childhood small noncleaved cell
C0281708|T191|Recurrent Childhood Burkitt's Lymphoma
C0281708|T191|Recurrent Pediatric Small Non-Cleaved Cell Lymphoma
C0281708|T191|childhood small noncleaved cell lymphoma, relapsed
C0281708|T191|Relapsed Pediatric Small Non-Cleaved Cell Lymphoma
C0281708|T191|Relapsed Childhood Small Non-Cleaved Cell Lymphoma
C0281708|T191|relapsed small noncleaved cell lymphoma, childhood
C0281708|T191|small noncleaved cell lymphoma, childhood, recurrent
C1956002|T045|Indel Mutation
C1956002|T045|Mutations, Insertion-Deletion
C1956002|T045|Insertion-Deletion Mutations
C1956002|T045|Mutations, INDEL
C1956002|T045|Insertion-Deletion Mutation
C1956002|T045|Mutation, Insertion-Deletion
C1956002|T045|Mutation, INDEL
C1956002|T045|Indel
C1956002|T045|INDEL Mutations
C1956002|T045|INDEL Mutation
C1956002|T045|Insertion Deletion Mutation
C1334160|T191|Immunodeficiency-Related Malignant Neoplasm
C1334160|T191|Immunosuppression-Related Malignant Neoplasm
C1334160|T191|Immunosuppression-Related Malignancy
C1334160|T191|Immunosuppression-Related Cancer
C0854798|T191|Recurrent Hepatoblastoma
C0854798|T191|Relapsed Hepatoblastoma
C0854798|T191|Hepatoblastoma, Recurrent
C0854798|T191|Hepatoblastoma recurrent
C0278649|T191|Recurrent Childhood Rhabdomyosarcoma
C0278649|T191|recurrent pediatric rhabdomyosarcoma
C0278649|T191|rhabdomyosarcoma, recurrent childhood
C0278649|T191|childhood rhabdomyosarcoma, recurrent
C0278649|T191|pediatric rhabdomyosarcoma, recurrent
C0278649|T191|Recurrent Pediatric Rhabdomyosarcoma
C0278649|T191|Relapsed Childhood Rhabdomyosarcoma
C0278649|T191|Relapsed Pediatric Rhabdomyosarcoma
C0278649|T191|recurrent childhood rhabdomyosarcoma
C1541273|T191|Recurrent Marginal Zone Lymphoma
C1541273|T191|recurrent marginal zone B-cell lymphoma
C1541273|T191|recurrent marginal zone lymphoma
C1541273|T191|Recurrent Marginal Zone B-Cell Lymphoma
C1335429|T191|Plasmacytoma-Like Post-Transplant Lymphoproliferative Disorder
C1335429|T191|Plasmacytoma-like PTLD
C3468050|T191|Adult Anaplastic (Malignant) Meningioma
C3468050|T191|Adult Anaplastic Meningioma
C3468050|T191|Adult Malignant Meningioma
C116542|T061|Pulsed-Dose Rate Brachytherapy
C0445064|T033|M1b Stage Finding
C0445064|T033|Metastasis stage M1b (finding)
C0445064|T033|M1b TNM Finding
C0445064|T033|Metastasis Stage M1b
C0445064|T033|M1b Distant Metastasis Stage Finding
C0445064|T033|Metastasis stage M1b
C0445064|T033|M1b Metastasis Finding
C0445064|T033|M1b Cancer Stage Finding
C0445064|T033|M1b
C0445064|T033|M1b Metastasis Stage
C0445064|T033|M1b Stage
C0445064|T033|M1b Distant Metastasis Finding
C1302494|T201|Size of base of tumor on transillumination, dimension 2
C1302494|T201|Size of base of tumour on transillumination, dimension 2
C1302494|T201|Size of base of tumor on transillumination, dimension 2 (observable entity)
C0279838|T191|Recurrent Oropharyngeal Carcinoma
C0279838|T191|recurrent carcinoma of the oropharynx
C0279838|T191|recurrent cancer of the oropharynx
C0279838|T191|Recurrent Oropharynx Carcinoma
C0279838|T191|oropharyngeal cancer, recurrent
C0279838|T191|Relapsed Cancer of the Oropharynx
C0279838|T191|recurrent oropharynx carcinoma
C0279838|T191|Relapsed Carcinoma of Oropharynx
C0279838|T191|Relapsed Cancer of Oropharynx
C0279838|T191|Relapsed Oropharynx Carcinoma
C0279838|T191|Recurrent Oropharyngeal Cancer
C0279838|T191|relapsed oropharyngeal carcinoma
C0279838|T191|Recurrent Cancer of Oropharynx
C0279838|T191|recurrent carcinoma of oropharynx
C0279838|T191|Recurrent Carcinoma of the Oropharynx
C0279838|T191|Relapsed Carcinoma of the Oropharynx
C0279838|T191|Oropharyngeal cancer recurrent
C0279838|T191|relapsed oropharyngeal cancer
C0279838|T191|Recurrent Cancer of the Oropharynx
C0279838|T191|relapsed cancer of the oropharynx
C0279838|T191|oropharynx cancer, recurrent
C0279838|T191|recurrent oropharyngeal cancer
C0279838|T191|relapsed carcinoma of the oropharynx
C0279838|T191|Relapsed Oropharyngeal Carcinoma
C0279838|T191|recurrent cancer of oropharynx
C0279838|T191|Oropharyngeal Cancer, Recurrent
C0279838|T191|Recurrent Carcinoma of Oropharynx
C0279838|T191|relapsed carcinoma of oropharynx
C0279838|T191|Relapsed Oropharyngeal Cancer
C0279838|T191|relapsed oropharynx carcinoma
C0279838|T191|relapsed cancer of oropharynx
C0441906|T033|V0 stage
C0441906|T033|V0 Stage
C0441906|T033|V0 Cancer Stage Finding
C0441906|T033|Venous Stage V0
C0441906|T033|V0 Stage Finding
C0441906|T033|V0
C0441906|T033|V0 Venous Invasion Finding
C0441906|T033|V0 Venous Stage
C0441906|T033|V0 stage (finding)
C0441906|T033|V0 TNM Finding
C0441906|T033|Venous stage V0
C0441906|T033|V0: no venous invasion
C0280097|T191|Squamous Cell Carcinoma of Unknown Primary Origin
C0280097|T191|Squamous Cell Carcinoma of Unknown Primary
C1335461|T191|Postsurgical Stage I Hepatoblastoma
C1302460|T201|Size of base of tumor on transillumination, dimension 1
C1302460|T201|Size of base of tumour on transillumination, dimension 1
C1302460|T201|Size of base of tumor on transillumination, dimension 1 (observable entity)
C2986683|T191|Stage I AIDS-Related Lymphoma
C2986683|T191|stage I AIDS-related lymphoma
C0346975|T191|Metastatic Malignant Neoplasm to the Rectum
C0346975|T191|Metastatic Tumor to the Rectum
C0346975|T191|Metastatic Neoplasm to the Rectum
C0346975|T191|Metastasis to the Rectum
C1332052|T191|AIDS-Related Non-Hodgkin Lymphoma of the Cervix
C1332052|T191|AIDS-Related Non-Hodgkin's Lymphoma of Cervix
C1332052|T191|AIDS-Related Non-Hodgkin's Lymphoma of the Cervix
C1332052|T191|AIDS-Related Uterine Cervical Non-Hodgkin's Lymphoma
C0854742|T191|Recurrent AIDS-Related Anal Canal Carcinoma
C0854742|T191|Recurrent AIDS-Related Anal Carcinoma
C0854742|T191|Recurrent AIDS-Related Anal Canal Cancer
C0854742|T191|Recurrent AIDS-Related Anal Cancer
C0278601|T191|Inflammatory Breast Carcinoma
C0278601|T191|Mastitis Carcinomatosa
C0278601|T191|carcinoma of the breast, inflammatory
C0278601|T191|Inflammatory Breast Neoplasms
C0278601|T191|Mastitis carcinomatosa
C0278601|T191|Inflammatory carcinoma of breast (disorder)
C0278601|T191|Inflammatory Breast Carcinomas
C0278601|T191|Inflammatory Breast Cancer
C0278601|T191|Inflammatory Breast Neoplasms [Disease/Finding]
C0278601|T191|Cancers, Inflammatory Breast
C0278601|T191|Inflammatory Breast Cancers
C0278601|T191|Neoplasm, Inflammatory Breast
C0278601|T191|Breast Carcinoma, Inflammatory
C0278601|T191|Cancer, Inflammatory Breast
C0278601|T191|Inflammatory Carcinoma of Breast
C0278601|T191|Inflammatory breast carcinoma
C0278601|T191|Inflammatory carcinoma of breast
C0278601|T191|Breast Carcinomas, Inflammatory
C0278601|T191|Inflammatory Breast Neoplasm
C0278601|T191|Breast Cancers, Inflammatory
C0278601|T191|Neoplasms, Inflammatory Breast
C0278601|T191|Inflammatory carcinoma of the breast
C0278601|T191|Carcinomas, Inflammatory Breast
C0278601|T191|Breast carcinoma inflammatory
C0278601|T191|Inflammatory breast cancer
C0278601|T191|Carcinoma, Inflammatory Breast
C0278601|T191|Inflammatory Breast Cancer (IBC)
C0278601|T191|inflammatory breast cancer
C0278601|T191|Breast Neoplasms, Inflammatory
C0278601|T191|Breast Neoplasm, Inflammatory
C0278601|T191|Breast Cancer, Inflammatory
C0278601|T191|Inflammatory Carcinoma of the Breast
C0278601|T191|breast cancer, inflammatory
C0279616|T191|Childhood Botryoid-Type Embryonal Rhabdomyosarcoma
C0279616|T191|Childhood Botryoid Rhabdomyosarcoma
C0279616|T191|Childhood Sarcoma Botryoides
C1514692|T061|Radiation Non-Ionizing, Radiotherapy
C1880036|T061|Chemotherapy Regimen Used to Treat Breast Carcinoma
C1518167|T191|Malignant Breast Myoepithelioma
C1518167|T191|Breast Myoepithelial Carcinoma
C1332976|T191|Childhood Leptomeningeal Melanoma
C1332976|T191|Pediatric Leptomeningeal Melanoma
C0424861|T033|Diameter of lump
C0424861|T033|Diameter of lump (observable entity)
C111695|T191|Mesenchymal Glioblastoma
C0424860|T033|Lump size
C0424860|T033|Size of mass
C0424860|T033|Lump size (observable entity)
C0424860|T033|Size of lump
C1711205|T033|Painless Mass
C0279019|T061|Mixed High-Low LET Therapy
C1515868|T191|Acinic Cell Breast Carcinoma
C1512908|T033|Intestinal Ulcerated Mass
C1879995|T061|Capecitabine-Docetaxel Regimen
C1879995|T061|XT Regimen
C1333285|T191|Diencephalic Glioblastoma
C1333285|T191|Grade IV Diencephalic Astrocytic Neoplasm
C1333285|T191|Grade IV Astrocytic Tumor of Diencephalon
C1333285|T191|Grade IV Astrocytic Neoplasm of the Diencephalon
C1333285|T191|Grade IV Astrocytic Neoplasm of Diencephalon
C1333285|T191|Glioblastoma Multiforme of Diencephalon
C1333285|T191|Diencephalic Glioblastoma Multiforme
C1333285|T191|GBM of the Diencephalon
C1333285|T191|Grade IV Diencephalic Astrocytic Tumor
C1333285|T191|Grade IV Astrocytic Tumor of the Diencephalon
C1333285|T191|Glioblastoma Multiforme of the Diencephalon
C1333285|T191|Diencephalic GBM
C1333285|T191|GBM of Diencephalon
C1333285|T191|Diencephalic Grade IV Astrocytoma
CL376151|T191|Childhood Favorable Prognosis Hodgkin Lymphoma
CL376151|T191|childhood favorable prognosis Hodgkin lymphoma
C2827415|T061|Radioactive Instillation
C0404186|T061|Right Salpingo-Oophorectomy
C1334743|T191|Metastatic Squamous Cell Breast Carcinoma
C1334743|T191|Metastatic Squamous Cell Carcinoma of the Breast
C1334743|T191|Metastatic Squamous Cell Carcinoma of Breast
C0686619|T191|Metastatic Malignant Neoplasm to the Lymph Node
C0686619|T191|Metastatic Tumor to Lymph Node
C0686619|T191|Metastatic Neoplasm to the Lymph Node
C0686619|T191|Metastasis to Lymph Node
C0686619|T191|Metastases to Lymph Nodes
C1519368|T191|Anaplastic Large Cell Lymphoma, Giant Cell Rich Subtype
C103267|T201|Narrow Surgical Margin
C103267|T201|Close Surgical Margin
C0279645|T191|Childhood Acute Monoblastic Leukemia
C0279645|T191|M5a leukemia, childhood acute
C0279645|T191|Childhood Acute M5a Leukemia
C0279645|T191|acute monocytic leukemia without differentiation, childhood
C0279645|T191|M5a Childhood Acute Monoblastic Leukemia without Differentiation
C0279645|T191|pediatric acute M5a leukemia
C0279645|T191|pediatric acute monocytic leukemia without differentiation
C0279645|T191|M5a childhood acute monocytic leukemia without differentiation
C0279645|T191|leukemia, childhood acute monocytic without differentiation
C0279645|T191|M5a childhood acute poorly differentiated monocytic leukemia
C0279645|T191|acute monoblastic leukemia, childhood
C0279645|T191|M5a Pediatric Acute Monoblastic Leukemia without Differentiation
C0279645|T191|pediatric acute poorly differentiated monocytic leukemia
C0279645|T191|leukemia, pediatric acute monoblastic
C0279645|T191|monoblastic leukemia, childhood acute
C0279645|T191|childhood acute monoblastic leukemia (M5a)
C0279645|T191|M5a pediatric acute monocytic leukemia without differentiation
C0279645|T191|Pediatric Acute Monoblastic Leukemia without Differentiation
C0279645|T191|pediatric AMOL, poorly differentiated
C0279645|T191|Pediatric Acute M5a Leukemia
C0279645|T191|Childhood Acute Monoblastic Leukemia without Differentiation
C0279645|T191|pediatric acute monoblastic leukemia
C0279645|T191|childhood acute poorly differentiated monocytic leukemia (M5a)
C0279645|T191|childhood acute monocytic leukemia without differentiation
C0279645|T191|childhood AMOL, poorly differentiated
C0279645|T191|childhood acute M5a leukemia
C2826148|T191|Therapy-Related Myelodysplastic/Myeloproliferative Neoplasm
C2826148|T191|Therapy-Related Myelodysplastic/Myeloproliferative Disease
C2826148|T191|t-MDS/MPN
C1515866|T191|Acinar Prostate Adenocarcinoma, Pseudohyperplastic Variant
C0279696|T191|Squamous Cell Carcinoma Metastatic to the Neck with Occult Primary
C0279696|T191|Metastatic Epidermoid Neck Cancer with Occult Primary
C0279696|T191|Metastatic Squamous Neck Cancer with Occult Primary
C0279696|T191|Squamous Cell Cancer Metastatic to the Neck with Occult Primary
C0279696|T191|Epidermoid Cancer Metastatic to the Neck with Occult Primary
C0279696|T191|Metastatic Squamous Cell Neck Cancer with Occult Primary
C0279696|T191|Squamous Cell Cancer Metastatic to Neck, with Occult Primary
C1709926|T170|Response Evaluation Criteria in Solid Tumors
C1709926|T170|RECIST
C1879500|T061|AC-T Regimen
C1879500|T061|AC-Taxol regimen
C1879500|T061|AC-T regimen
C1879500|T061|AC-Taxol Regimen
C1879500|T061|AC-T
C0454271|T061|Low-Dose Rate Brachytherapy
C1332233|T191|Alkylating Agent-Related Acute Myeloid Leukemia
C1332233|T191|Alkylating Agent-Related AML
C1332233|T191|Alkylating Agent Related Acute Myeloid Leukemia
C1706789|T191|Ameloblastic Carcinoma-Secondary Type (Dedifferentiated), Intraosseous
C1706789|T191|Central Ameloblastic Carcinoma
C2348909|T034|HER2/Neu Positive
C2348909|T034|ERBB2 Positive
C111241|T061|Laser Ablation
C111241|T061|Ablation, Laser
C111241|T061|Laser Tissue Ablation
C111241|T061|Laser Photoablation of Tissue
C111241|T061|Vaporization, Laser
C111241|T061|Vaporization
C111241|T061|Tissue Ablation, Laser
C111241|T061|Photoablation
C111241|T061|Ablation, Laser Tissue
C111241|T061|Laser ablation
C111241|T061|Laser Vaporization
C111241|T061|Pulsed Laser Tissue Ablation
C111241|T061|ABLATION, LASER
C2919529|T081|Calculated volume of neoplasm using magnetic resonance imaging
C2919529|T081|Calculated volume of neoplasm using magnetic resonance imaging (observable entity)
C0475413|T033|Tumor stage Tis
C0475413|T033|Tis Stage Finding
C0475413|T033|Tis Tumor Finding
C0475413|T033|Tis TNM Finding
C0475413|T033|Tis category (finding)
C0475413|T033|Tis: Carcinoma in situ
C0475413|T033|Tis Cancer Stage Finding
C0475413|T033|Tis Stage
C0475413|T033|Tis Tumor Stage
C0475413|T033|Tis Primary Tumor Stage Finding
C0475413|T033|Tis category
C0475413|T033|Tis stage
C0475413|T033|Tis
C0475413|T033|Tumour stage Tis
C0475413|T033|Tis Primary Tumor Finding
C0475413|T033|Tumor Stage Tis
C0220654|T191|Meningeal Carcinomatosis
C0220654|T191|Meningeal carcinomatosis
C0220654|T191|Lymphomatous meningitis
C0220654|T191|INTRACRANIAL NEOPLASM, MENINGEAL CARCINOMATOSIS
C0220654|T191|neoplastic meningitis
C0220654|T191|Meningitis, Carcinomatous
C0220654|T191|Carcinomatosis of the Meninges
C0220654|T191|carcinomatous leptomeningitis
C0220654|T191|meningitis, carcinomatous
C0220654|T191|Carcinomatous Meningitides
C0220654|T191|MENINGEAL CARCINOMATOSIS
C0220654|T191|Leptomeningeal Carcinomatoses
C0220654|T191|BRAIN TUMOR, MENINGEAL CARCINOMATOSIS
C0220654|T191|Carcinomatosis, Leptomeningeal
C0220654|T191|Leptomeningeal Carcinomatosis
C0220654|T191|Carcinomatoses, Leptomeningeal
C0220654|T191|Meningeal Carcinomatoses
C0220654|T191|Malignant meningitis (disorder)
C0220654|T191|meningeal carcinomatosis
C0220654|T191|Meningeal Carcinomatosis [Disease/Finding]
C0220654|T191|Neoplastic meningitis
C0220654|T191|Meningitides, Carcinomatous
C0220654|T191|CANCER, MENINGEAL CARCINOMATOSIS
C0220654|T191|carcinomatous meningitis
C0220654|T191|Carcinomatosis, Meningeal
C0220654|T191|Carcinomatoses, Meningeal
C0220654|T191|Carcinomatous Meningitis
C0220654|T191|Carcinomatous meningitis
C0220654|T191|Malignant meningitis
C0476661|T033|Prophylactic Surgery
C0476661|T033|Prophylactic surgery, unspecified
C0476661|T033|Prophylactic surgery
C0476661|T033|prophylactic surgery
C0476661|T033|Encounter due to prophylactic surgery, unspecified
C0854777|T191|Recurrent Pancreatic Carcinoma
C0854777|T191|Relapsed Cancer of the Pancreas
C0854777|T191|Recurrent Pancreatic Cancer
C0854777|T191|Recurrent Carcinoma of the Pancreas
C0854777|T191|Pancreatic carcinoma recurrent
C0854777|T191|recurrent pancreatic cancer
C0854777|T191|Pancreatic Carcinoma, Recurrent
C0854777|T191|Relapsed Pancreatic Carcinoma
C0854777|T191|pancreas cancer, recurrent
C0854777|T191|Recurrent Cancer of the Pancreas
C0854777|T191|recurrent pancreas cancer
C0854777|T191|Pancreas carcinoma recurrent
C0854777|T191|Relapsed Pancreatic Cancer
C0854777|T191|Pancreatic cancer recurrent
C0854777|T191|Recurrent Carcinoma of Pancreas
C0854777|T191|Relapsed Carcinoma of the Pancreas
C0854777|T191|Relapsed Cancer of Pancreas
C0854777|T191|pancreatic cancer, recurrent
C0854777|T191|Recurrent Cancer of Pancreas
C0854777|T191|Relapsed Carcinoma of Pancreas
C1332943|T191|Childhood Anaplastic Oligodendroglioma
C1332943|T191|anaplastic childhood oligodendroglioma
C1332943|T191|Anaplastic Childhood Oligodendroglioma
C1332943|T191|anaplastic pediatric oligodendroglioma
C1332943|T191|Undifferentiated Childhood Oligodendroglioma
C1332943|T191|childhood anaplastic oligodendroglioma
C1332943|T191|Undifferentiated Pediatric Oligodendroglioma
C1332943|T191|undifferentiated pediatric oligodendroglioma
C1332943|T191|Anaplastic Pediatric Oligodendroglioma
C1332943|T191|undifferentiated childhood oligodendroglioma
C0334246|T191|Metastatic Squamous Cell Carcinoma
C0334246|T191|Metastatic squamous cell carcinoma (disorder)
C0334246|T191|Squamous cell carcinoma, metastatic
C0334246|T191|Squamous cell carcinoma, metastatic, NOS
C0334246|T191|Squamous cell carcinoma, metastatic (morphologic abnormality)
C0334246|T191|Metastatic squamous cell carcinoma
C0278623|T061|High-LET Neutron Therapy
C0278623|T061|fast-neutron beam radiation
C0278623|T061|therapy, neutron
C0278623|T061|therapy, high-LET neutron
C0278623|T061|neutron therapy
C1336813|T191|Transplant-Related Lung Carcinoma
C1321214|T033|Tumor size, left ovary
C1321214|T033|Tumour size, left ovary
C1321214|T033|Tumor size, left ovary (observable entity)
C1708656|T191|Laryngeal Squamous Cell Carcinoma, Spindle Cell Variant
C1708656|T191|Laryngeal Carcinosarcoma
C1708656|T191|Laryngeal Sarcomatoid Carcinoma
C1512419|T191|Hereditary Melanoma
C1512419|T191|Melanoma, Familial
C1512419|T191|melanoma, hereditary, multiple
C1512419|T191|Hereditary Cutaneous Melanoma
C1512419|T191|Familial Melanoma
C1512419|T191|hereditary multiple melanoma
C1512419|T191|Familial Cutaneous Melanoma
C0850292|T061|Radiofrequency Ablation
C0850292|T061|Radiofrequency Interstitial Ablation
C0850292|T061|radiofrequency ablation
C0850292|T061|Radiofrequency ablation
C0279982|T191|Childhood Synovial Sarcoma
C0279982|T191|pediatric synovial sarcoma
C0279982|T191|Pediatric Synovial Sarcoma
C0279982|T191|sarcoma, synovial, childhood
C0279982|T191|synovial sarcoma, childhood
C0279982|T191|childhood synovial sarcoma
C0279982|T191|synovial sarcoma, pediatric
C2985448|T191|Radiation-Related Sarcoma
C3273930|T033|Tumor Mass
C3273930|T033|Tumor
C1512740|T191|Infiltrating Bladder Urothelial Carcinoma, Microcystic Variant
C0563529|T061|Left Oophorectomy
C0563529|T061|Left oophorectomy (procedure)
C0563529|T061|Left oophorectomy
C0563529|T061|Oophorectomy left
C0475395|T185|T4a Stage Finding
C0475395|T185|T4a Primary Tumor Finding
C0475395|T185|T4a
C0475395|T185|T4a Stage
C0475395|T185|Tumour stage T4a
C0475395|T185|T4a Tumor Finding
C0475395|T185|Tumor Stage T4a
C0475395|T185|T4a TNM Finding
C0475395|T185|Tumor stage T4a
C0475395|T185|T4a Tumor Stage
C0475395|T185|T4a Cancer Stage Finding
C0475395|T185|T4a tumor stage
C0475395|T185|T4a Primary Tumor Stage Finding
C0475395|T185|Tumor stage T4a (finding)
C1142163|T047|Intestinal Mass
C1142163|T047|Intestinal mass
C1335983|T191|Small Cell Variant Anaplastic Large Cell Lymphoma
C0278556|T191|Recurrent Anal Canal Carcinoma
C0278556|T191|recurrent anus cancer
C0278556|T191|recurrent anal cancer
C0278556|T191|Recurrent Anal Cancer
C0278556|T191|anus cancer, recurrent
C0278556|T191|Anal carcinoma recurrent
C0278556|T191|Anal canal cancer recurrent
C0278556|T191|anal cancer, recurrent
C0278556|T191|Anal cancer recurrent
C0278556|T191|Recurrent Anal Canal Cancer
C0854851|T191|Recurrent Mature T- and NK-Cell Non-Hodgkin Lymphoma
C0854851|T191|Relapsed Peripheral T-cell Lymphoma
C0854851|T191|Recurrent Peripheral T-cell Lymphoma
C0854851|T191|Recurrent Mature T- and NK-Cell Lymphoma
C0854851|T191|Recurrent Mature T- and NK-Cell Non-Hodgkin's Lymphoma
C1336023|T191|Solar Radiation-Related Skin Melanoma
C1336023|T191|Solar Radiation-Related Melanoma of the Skin
C1336023|T191|Solar Radiation-Related Melanoma of Skin
CL018755|T191|Ductal Breast Carcinoma In Situ and Invasive Lobular Carcinoma
CL018755|T191|DCIS and Infiltrating Lobular Carcinoma
CL018755|T191|Non-Infiltrating Ductal Carcinoma and ILC
CL018755|T191|DCIS and ILC
CL018755|T191|Non-Infiltrating Ductal Carcinoma and Infiltrating Lobular Carcinoma
CL018755|T191|Ductal Carcinoma in situ and Infiltrating Lobular Carcinoma
C1541469|T191|Recurrent Adult Grade III Lymphomatoid Granulomatosis
C1336812|T191|Transplant-Related Kaposi Sarcoma
C1336812|T191|Transplant-Related Kaposi's Sarcoma
C0278512|T191|Metastatic Osteosarcoma
C0278512|T191|sarcoma, metastatic osteogenic
C0278512|T191|metastatic osteosarcoma
C0278512|T191|metastatic osteogenic sarcoma
C0278512|T191|osteogenic sarcoma, metastatic
C0278512|T191|Metastatic Osteogenic Sarcoma
C0278512|T191|Osteosarcoma metastatic
C0278512|T191|Osteosarcoma, Metastatic
C0278512|T191|osteosarcoma, metastatic
C0278512|T191|Osteogenic sarcoma metastatic
C0854821|T191|Refractory Anaplastic Large Cell Lymphoma
C0854821|T191|Anaplastic Large Cell Lymphoma T- and Null-cell Types Refractory
C0854821|T191|Anaplastic large cell lymphoma T- and null-cell types refractory
CL388429|T191|Childhood Anaplastic Oligoastrocytoma
CL388429|T191|childhood oligoastrocytoma
CL388429|T191|childhood gliomas, mixed
CL388429|T191|childhood tumors, mixed glial
CL388429|T191|childhood mixed glioma
CL388429|T191|Brain tumor, child: Mixed glioma
CL388429|T191|childhood anaplastic oligoastrocytoma
CL388429|T191|childhood mixed glial tumors
CL388429|T191|childhood glial tumors, mixed
CL388429|T191|Childhood Mixed Glioma
C1335426|T191|Plasma Cell Post-Transplant Lymphoproliferative Disorder
C1335426|T191|Plasma Cell PTLD
C1704231|T191|Secondary Central Nervous System Lymphoma
C1704231|T191|meningitis, lymphomatous
C1704231|T191|Lymphomatous meningitis (disorder)
C1704231|T191|lymphomatous leptomeningitis
C1704231|T191|Lymphomatous meningitis
C1704231|T191|lymphomatous meningitis
C1704231|T191|secondary central nervous system lymphoma
C1704231|T191|leptomeningitis, lymphomatous
C1332059|T191|AIDS-Related Primary Effusion Lymphoma
C1301092|T201|Maximal height of tumor, after sectioning
C1301092|T201|Maximal height of tumor, after sectioning (observable entity)
C1301092|T201|Maximal height of tumour, after sectioning
C2348910|T034|HER2/Neu Status Unknown
C115292|T191|Non-Metastatic Childhood Soft Tissue Sarcoma
C3273076|T191|Extrarenal Rhabdoid Tumor of the Liver
C3273076|T191|Extrarenal Malignant Rhabdoid Tumor of the Liver
C2985561|T061|Total Skin Electron Beam Radiation Therapy
C2985561|T061|total skin electron beam radiation therapy
C2985561|T061|TSEB radiation therapy
C1334216|T191|Intermediate Grade Malignant Neoplasm
C1879523|T061|AT Regimen
C1879523|T061|Adriamycin-Taxol Regimen
C0279983|T191|Malignant Childhood Hemangiopericytoma
C0279983|T191|hemangiopericytoma, malignant, childhood
C0279983|T191|childhood malignant hemangiopericytoma
C0279983|T191|Childhood Malignant Hemangiopericytoma
C0279983|T191|Malignant Pediatric Hemangiopericytoma
C0279983|T191|malignant hemangiopericytoma, pediatric
C0279983|T191|malignant hemangiopericytoma, childhood
C0279983|T191|pediatric malignant hemangiopericytoma
C1519182|T191|Skin Sarcomatoid Basal Cell Carcinoma
C0475374|T033|T3 Stage Finding
C0475374|T033|T3 stage
C0475374|T033|T3 TNM Finding
C0475374|T033|T3 category (finding)
C0475374|T033|Tumor Stage T3
C0475374|T033|T3 category
C0475374|T033|T3 Tumor Stage
C0475374|T033|T3 Primary Tumor Finding
C0475374|T033|T3 Cancer Stage Finding
C0475374|T033|T3
C0475374|T033|Tumour stage T3
C0475374|T033|T3 Primary Tumor Stage Finding
C0475374|T033|Tumor stage T3
C0475374|T033|T3 Stage
C0475374|T033|T3 tumor stage
C0475374|T033|T3 Tumor Finding
C1334407|T191|Localized Carcinoma
C1334407|T191|Localized Cancer
C1332549|T191|Bilateral Carcinoma
C1332549|T191|Bilateral Cancer
C1332549|T191|bilateral cancer
C0862641|T191|Stage II Prostate Adenocarcinoma
C0862641|T191|Stage II Prostate Adenocarcinoma AJCC v7
C1708232|T033|Generic Regional Lymph Nodes TNM Finding
C0854793|T191|Non-Resectable Malignant Liver Neoplasm
C0854793|T191|Non-Resectable Hepatic Malignant Neoplasm
C0854793|T191|Non-Resectable Malignant Neoplasm of Liver
C1710523|T049|UV Mutation Abnormality
C1710523|T049|UV-Mutagenesis
C2985559|T061|Plaque Radiotherapy
C2985559|T061|plaque radiotherapy
C1332282|T191|Anaplastic Hemispheric Astrocytoma
C1332282|T191|Grade III Astrocytic Tumor of Cerebral Hemisphere
C1332282|T191|Anaplastic Astrocytoma of Cerebral Hemisphere
C1332282|T191|Anaplastic Astrocytoma, Hemispheric
C1332282|T191|Grade III Cerebral Hemisphere Astrocytic Neoplasm
C1332282|T191|Grade III Cerebral Hemisphere Astrocytic Tumor
C1332282|T191|Grade III Astrocytoma of Cerebral Hemisphere
C1332282|T191|Anaplastic Astrocytoma of the Cerebral Hemisphere
C1332282|T191|Grade III Hemispheric Astrocytic Neoplasm
C1332282|T191|Grade III Astrocytic Neoplasm of Cerebral Hemisphere
C1332282|T191|Grade III Hemispheric Astrocytic Tumor
C1332282|T191|Undifferentiated Astrocytoma of the Cerebral Hemisphere
C1332282|T191|Grade III Astrocytic Neoplasm of the Cerebral Hemisphere
C1332282|T191|Cerebral Hemisphere Anaplastic Astrocytoma
C1332282|T191|Grade III Cerebral Hemisphere Astrocytoma
C1332282|T191|Grade III Astrocytoma of the Cerebral Hemisphere
C1332282|T191|Hemispheric Anaplastic Astrocytoma
C1332282|T191|Undifferentiated Astrocytoma of Cerebral Hemisphere
C1332282|T191|Grade III Hemispheric Astrocytoma
C1332282|T191|Grade III Astrocytic Tumor of the Cerebral Hemisphere
C1335712|T191|Recurrent Medulloblastoma
C1335712|T191|Relapsed Medulloblastoma
C1335712|T191|Medulloblastoma recurrent
C1881206|T045|Inframe Mutation
C1335502|T191|Prostate Adenoid Cystic Carcinoma
C1335502|T191|Adenoid Cystic Carcinoma of Prostate
C1335502|T191|Adenoid Cystic Carcinoma of the Prostate
C0006413|T191|Childhood Burkitt Lymphoma
C0006413|T191|childhood small non-cleaved cell lymphoma
C0006413|T191|Burkitts Lymphoma
C0006413|T191|Burkitt's tumour or lymphoma
C0006413|T191|Pediatric Small Non-Cleaved Cell Lymphoma
C0006413|T191|Burkitt's tumour [obs]
C0006413|T191|LYMPHOMA, BURKITT
C0006413|T191|Leukemia, Burkitt's
C0006413|T191|Burkitt's tumor non-Hodgkin's lymphoma
C0006413|T191|Pediatric Burkitt's Lymphoma
C0006413|T191|BL - Burkitt's lymphoma
C0006413|T191|Burkitt Tumor
C0006413|T191|[M]Burkitt's tumour
C0006413|T191|Burkitt's lymphoma (clinical)
C0006413|T191|Burkitt Cell Leukemia
C0006413|T191|diffuse undifferentiated lymphoma, childhood
C0006413|T191|Childhood Small Non-Cleaved Cell Lymphoma
C0006413|T191|Leukemia, Lymphocytic, L3
C0006413|T191|Tumor, Burkitt's
C0006413|T191|lymphoma, Burkitt's
C0006413|T191|Burkitt Leukemia
C0006413|T191|Burkitt lymphoma (morphologic abnormality)
C0006413|T191|small noncleaved cell lymphoma, childhood
C0006413|T191|Leukemias, L3 Lymphocytic
C0006413|T191|Burkitt's lymphoma (disorder)
C0006413|T191|lymphoma, small non-cleaved cell, childhood
C0006413|T191|Leukemia, Burkitt
C0006413|T191|Burkitt's Leukemia
C0006413|T191|Burkitt lymphoma
C0006413|T191|Burkitt's type malignant lymphoma - small non-cleaved
C0006413|T191|NHL, Burkitt's
C0006413|T191|pediatric small non-cleaved cell lymphoma
C0006413|T191|childhood SNC lymphoma
C0006413|T191|Leukemia, Lymphoblastic, Burkitt-Type
C0006413|T191|childhood small noncleaved cell lymphoma
C0006413|T191|pediatric SNC lymphoma
C0006413|T191|Lymphoma, Burkitt
C0006413|T191|Malignant lymphoma, small noncleaved, Burkitt type [obs]
C0006413|T191|Small Non-Cleaved Cell Lymphoma, Burkitt's Type
C0006413|T191|lymphoma, small noncleaved cell, childhood
C0006413|T191|Burkitt tumor [obs]
C0006413|T191|DUL, childhood
C0006413|T191|Lymphocytic Leukemias, L3
C0006413|T191|Burkitt's lymphoma
C0006413|T191|Burkitt lymphoma, unspecified site
C0006413|T191|L3 Lymphocytic Leukemias
C0006413|T191|SNC lymphoma, childhood
C0006413|T191|small non-cleaved cell lymphoma, childhood
C0006413|T191|Lymphoma, Burkitt's
C0006413|T191|Burkitt's tumor [obs]
C0006413|T191|Burkitt's Lymphoma
C0006413|T191|Malignant lymphoma, Burkitt's type
C0006413|T191|Burkitt's lymphoma - disorder
C0006413|T191|Burkitt's tumor
C0006413|T191|Burkitt's type malignant lymphoma - undifferentiated
C0006413|T191|Burkitt Lymphoma
C0006413|T191|L3 Lymphocytic Leukemia
C0006413|T191|Burkitt's lymphomas
C0006413|T191|lymphoma, diffuse undifferentiated, childhood
C0006413|T191|BURKITT LYMPHOMA
C0006413|T191|Leukemia, Burkitt Cell
C0006413|T191|[M]Burkitt's tumor
C0006413|T191|Burkitt tumour [obs]
C0006413|T191|Burkitt's Tumor
C0006413|T191|BL
C0006413|T191|Lymphocytic Leukemia, L3
C0006413|T191|Malignant lymphoma, undifferentiated, Burkitt type [obs]
C0006413|T191|childhood Burkitt lymphoma
C0006413|T191|Burkitt's tumour
C0006413|T191|pediatric Burkitt lymphoma
C0006413|T191|Leukemia, L3 Lymphocytic
C0006413|T191|Burkitts Tumor
C0006413|T191|Tumor, Burkitt
C0006413|T191|Burkitt's lymphoma NOS
C0006413|T191|Burkitt's tumor or lymphoma
C0006413|T191|Malignant lymphoma, small noncleaved, Burkitt's, diffuse
C0006413|T191|Burkitts Leukemia
C0006413|T191|Burkitt lymphoma, NOS Includes all variants
C0006413|T191|Cell Leukemia, Burkitt
C0006413|T191|non-Hodgkin's lymphoma, Burkitt's
C0006413|T191|Childhood Burkitt's Lymphoma
C0006413|T191|Burkitt Lymphoma [Disease/Finding]
C1512745|T191|Infiltrating Bladder Urothelial Carcinoma, Sarcomatoid Variant without Heterologous Elements
C0279941|T191|Primary Childhood Soft Tissue Sarcoma
C0279941|T191|pediatric nonmetastatic STS
C0279941|T191|Nonmetastatic Childhood Soft Tissue Sarcoma
C0279941|T191|childhood STS, nonmetastatic
C0279941|T191|nonmetastatic childhood soft tissue sarcoma
C0279941|T191|Non-Metastatic Pediatric Soft Tissue Sarcoma
C0279941|T191|childhood soft tissue sarcoma, nonmetastatic
C0279941|T191|soft tissue sarcoma, nonmetastatic, childhood,
C0279941|T191|STS, nonmetastatic, childhood
C0279941|T191|Non-Metastatic Childhood Soft Tissue Sarcoma
C0279941|T191|childhood nonmetastatic STS
C0279941|T191|STS, childhood, nonmetastatic
C0279941|T191|pediatric STS, nonmetastatic
C0346158|T191|Juvenile Fibroadenoma
C0346158|T191|Cellular fibroadenoma
C0346158|T191|Juvenile fibroadenoma of breast (disorder)
C0346158|T191|Juvenile Breast Fibroadenoma
C0346158|T191|Juvenile fibroadenoma
C0346158|T191|Juvenile Fibroadenoma of Breast
C0346158|T191|Cellular Fibroadenoma
C0346158|T191|Juvenile Fibroadenoma of the Breast
C0346158|T191|Juvenile fibroadenoma of breast
C0346158|T191|Juvenile fibroadenoma (morphologic abnormality)
CL433909|T191|Childhood Giant Cell Glioblastoma
CL433909|T191|childhood giant cell glioblastoma
C0475386|T185|T1c Stage Finding
C0475386|T185|Tumor Stage T1c
C0475386|T185|T1c Cancer Stage Finding
C0475386|T185|T1c Primary Tumor Stage Finding
C0475386|T185|Tumour stage T1c
C0475386|T185|T1c Primary Tumor Finding
C0475386|T185|T1c Tumor Finding
C0475386|T185|T1c Stage
C0475386|T185|Tumor stage T1c (finding)
C0475386|T185|Tumor stage T1c
C0475386|T185|T1c
C0475386|T185|T1c Tumor Stage
C0475386|T185|T1c TNM Finding
C0449458|T082|Corticotroph adenoma size
C0449458|T082|Corticotroph adenoma size (observable entity)
C0449458|T082|Size of corticotroph adenoma
C0861819|T191|Metastatic Small Intestinal Adenocarcinoma
C0861819|T191|Small intestine adenocarcinoma metastatic
C0861819|T191|Small intestine adenocarcinoma metastatic NOS
C0855147|T191|Recurrent B Lymphoblastic Lymphoma
C0855147|T191|Recurrent B-Lymphoblastic Lymphoma
C0855147|T191|Relapsed Precursor B-Lymphoblastic Lymphoma
C0855147|T191|Recurrent Precursor B-Lymphoblastic Lymphoma
C0935764|T061|MRI-Guided Focused Ultrasound Ablation
C1377605|T191|Childhood Central Nervous System Embryonal Carcinoma
C1377605|T191|Embryonal Carcinoma of the Pediatric Central Nervous System
C1377605|T191|Embryonal Carcinoma of the Childhood Central Nervous System
C1377605|T191|Embryonal Carcinoma of the Childhood CNS
C1377605|T191|Embryonal Carcinoma of Childhood CNS
C1377605|T191|Embryonal Carcinoma of the Pediatric CNS
C1377605|T191|Embryonal Carcinoma of Pediatric Central Nervous System
C1377605|T191|Pediatric Central Nervous System Embryonal Carcinoma
C1377605|T191|Embryonal Carcinoma of Pediatric CNS
C1377605|T191|Embryonal Carcinoma of Childhood Central Nervous System
C1377605|T191|Pediatric CNS Embryonal Cell Carcinoma
C1377605|T191|Childhood CNS Embryonal Cell Carcinoma
CL448380|T191|Recurrent Carcinoma
CL448380|T191|Relapsed Cancer
CL448380|T191|Relapsed Carcinoma
CL448380|T191|Recurrent Cancer
C0919390|T121|Tamoxifen Citrate
C0919390|T121|Nolgen
C0919390|T121|Lesporene
C0919390|T121|Clonoxifen
C0919390|T121|(Z)-2-[4-(1,2-Diphenyl-1-butenyl)phenoxy]-N,N-dimethylethanamine 2-Hydroxy-1,2,3-propanetricarboxylate
C0919390|T121|Tamifen
C0919390|T121|(Z)-2-[4-(1,2-diphenyl-1-butenyl)phenoxy]-N,N-dimethylethanamine citrate
C0919390|T121|Nolvadex-D
C0919390|T121|Estroxyn
C0919390|T121|Emblon
C0919390|T121|tamoxifen citrate
C0919390|T121|Oestrifen
C0919390|T121|Tamaxin
C0919390|T121|Novofen
C0919390|T121|1-p-beta-dimethylamino-ethoxyphenyl-trans-1,2-diphenylbut-1-ene Citrate
C0919390|T121|Noxitem
C0919390|T121|TAM
C0919390|T121|Fentamox
C0919390|T121|Oncotam
C0919390|T121|Tamofen
C0919390|T121|TAMOXIFEN CITRATE
C0919390|T121|Kessar
C0919390|T121|Genox
C0919390|T121|Gen-Tamoxifen
C0919390|T121|Jenoxifen
C0919390|T121|Zemide
C0919390|T121|Apo-Tamox
C0919390|T121|Nolvadex
C0919390|T121|ICI 46,474
C0919390|T121|Ledertam
C0919390|T121|Tamax
C0919390|T121|Noltam
C0919390|T121|Tamoxifen citrate
C0919390|T121|Ebefen
C0919390|T121|Novo-Tamoxifen
C0919390|T121|Nourytam
C0919390|T121|Soltamox
C0919390|T121|PMS-Tamoxifen
C0919390|T121|Tamizam
C0919390|T121|Tamoxifeni Citras
C0919390|T121|Tamoxasta
C0919390|T121|ICI-46474
C0919390|T121|Dignotamoxi
C114950|T191|Secondary Central Nervous System Non-Hodgkin Lymphoma
C0278839|T191|Recurrent Skin Carcinoma
C0278839|T191|cancer of the skin, recurrent
C0278839|T191|skin cancer, recurrent
C0278839|T191|Recurrent Cancer of Skin
C0278839|T191|Recurrent Carcinoma of the Skin
C0278839|T191|recurrent skin cancer
C0278839|T191|Recurrent Cancer of the Skin
C0278839|T191|Recurrent Carcinoma of Skin
C0278839|T191|recurrent cancer of the skin
C0278839|T191|recurrent carcinoma of the skin
C0278839|T191|Recurrent Skin Cancer
C0278839|T191|Recurrent Cutaneous Carcinoma
C0278839|T191|carcinoma of the skin, recurrent
C1512814|T061|Intensity-Modulated Radiation Therapy
C1512814|T061|intensity-modulated radiation therapy
C1512814|T061|Intensity-Modulated Radiotherapy
C1512814|T061|IMRT
C1512814|T061|Intensity Modulated RT
C1512796|T045|Insertion Mutation
C1512796|T045|Mutations, Insertion
C1512796|T045|Insertion Mutation Abnormality
C1512796|T045|Insertion
C1512796|T045|Insertion Mutations
C1512796|T045|Mutation, Insertion
C0017086|T047|Gangrene
C0017086|T047|Gangrene [Disease/Finding]
C0017086|T047|Gangrenes
C0017086|T047|Gangrene, NOS
C0017086|T047|Gangrene ICD9CM:785.4
C0017086|T047|Gangrenous
C0017086|T047|Gangrene (morphologic abnormality)
C0017086|T047|Gangrenous disorder (disorder)
C0017086|T047|Gangrene NOS
C0017086|T047|gangrene
C0017086|T047|Gangrenous disorder
C0017086|T047|GANGRENE
C0445085|T033|NX Stage Finding
C0445085|T033|Node stage NX
C0445085|T033|NX
C0445085|T033|NX category (finding)
C0445085|T033|NX Lymph Node Stage
C0445085|T033|NX Lymph Node Finding
C0445085|T033|NX Stage
C0445085|T033|NX stage
C0445085|T033|NX Regional Lymph Nodes Finding
C0445085|T033|NX Cancer Stage Finding
C0445085|T033|Lymph Node Stage NX
C0445085|T033|NX Node Stage
C0445085|T033|NX category
C0445085|T033|NX Node Finding
C0445085|T033|NX TNM Finding
C0445085|T033|NX lymph node stage
C0445085|T033|NX Regional Lymph Node Stage Finding
C0445085|T033|Node Stage NX
C1265603|T190|Firm Mass
C1265603|T190|Firm mass
C1265603|T190|Firm mass (morphologic abnormality)
C0876982|T191|Unresectable Gallbladder Carcinoma
C0876982|T191|unresectable gallbladder cancer
C0876982|T191|gallbladder cancer, unresectable
C0876982|T191|Unresectable Gallbladder Cancer
C0876982|T191|Gallbladder Carcinoma Unresectable
C0876982|T191|Unresectable Cancer of Gallbladder
C0876982|T191|Gallbladder carcinoma non-resectable
C0876982|T191|Gallbladder Cancer Unresectable
C0876982|T191|Unresectable Cancer of the Gallbladder
C0876982|T191|Gallbladder cancer non-resectable
C1334275|T191|Invasive Cribriform Breast Carcinoma
C1334275|T191|Invasive Cribriform Carcinoma of Breast
C1334275|T191|Invasive Cribriform Carcinoma of the Breast
C1334275|T191|Infiltrating Cribriform Carcinoma of Breast
C1334275|T191|Infiltrating Cribriform Carcinoma of the Breast
C1334275|T191|Infiltrating Cribriform Breast Carcinoma
C1334275|T191|Infiltrating Cribriform Ductal Carcinoma of Breast
C1334275|T191|Invasive Cribriform Ductal Carcinoma of Breast
C0278884|T191|Recurrent Melanoma
C0278884|T191|Recurrent Malignant Melanoma
C0278884|T191|Melanoma recurrent
C0278884|T191|recurrent melanoma
C0278884|T191|melanoma, recurrent
C1332049|T191|AIDS-Related Malignant Anal Neoplasm
C1332049|T191|AIDS-Related Malignant Neoplasm of the Anus
C1332049|T191|AIDS-Related Malignant Tumor of the Anus
C1332049|T191|AIDS-Related Malignant Anal Tumor
C1332049|T191|AIDS-Related Malignant Neoplasm of Anus
C1332049|T191|AIDS-Related Malignant Tumor of Anus
C1879492|T061|A-CMF Regimen
C1879492|T061|Adriamycin-Cytoxan-Methotrexate-Fluorouracil Regimen
C1335752|T191|Infiltrating Renal Pelvis Urothelial Carcinoma, Sarcomatoid Variant
C1335752|T191|Sarcomatoid Transitional Cell Carcinoma of Renal Pelvis
C1335752|T191|Sarcomatoid Transitional Cell Carcinoma of the Renal Pelvis
C1335752|T191|Sarcomatoid Transitional Cell Carcinoma of Kidney Pelvis
C1335752|T191|Sarcomatoid Transitional Cell Carcinoma of the Kidney Pelvis
C1335752|T191|Kidney Pelvis Sarcomatoid Transitional Cell Carcinoma
C2987250|T191|Second Primary Malignant Neoplasm
C2987250|T191|Second Primary Cancer
C2987250|T191|second cancer
CL448482|T191|Recurrent Askin Tumor
CL448482|T191|Recurrent Askin's Tumor
C1403582|T081|Mass
C1403582|T081|Lung mass (finding)
C1403582|T081|BREAST MASS
C1403582|T081|Breast Lump
C1403582|T081|Lung Mass
C1403582|T081|subcutaneous mass
C1403582|T081|cutaneous mass
C1403582|T081|Breast Mass
C1403582|T081|MASS
C1403582|T081|Hepatic mass
C1403582|T081|Breast Nodule
C1403582|T081|area of enhancement
C1403582|T081|lesion
C1403582|T081|nodule
C1403582|T081|mass
C1403582|T081|SUBCUTANEOUS MASS
C1403582|T081|liver mass
C1403582|T081|Localized mass
C1403582|T081|molecular weight
C1403582|T081|Lumpy breast
C1403582|T081|Pulmonary mass
C1403582|T081|MOL WEIGHT
C1403582|T081|vague density
C1403582|T081|Mass (morphologic abnormality)
C1403582|T081|Mass (quantity of matter)
C1403582|T081|Breast mass NOS
C1403582|T081|Breast mass
C1403582|T081|Dermatologic Mass
C1403582|T081|Mass in Breast
C1403582|T081|epidermal mass
C1403582|T081|Mass, a measure of quantity of matter (property)
C1403582|T081|Mass, a measure of quantity of matter (property) (qualifier value)
C1403582|T081|mw
C1403582|T081|dermal mass
C1403582|T081|Lump or mass in breast
C1403582|T081|Mass of body structure (finding)
C1403582|T081|LUMPS, BREAST
C1403582|T081|focus
C1403582|T081|dermatologic mass
C1403582|T081|Molecular Weight
C1403582|T081|Weights, Molecular
C1403582|T081|Lung mass
C1403582|T081|Mass in breast
C1403582|T081|Mass NOS
C1403582|T081|Unspecified lump in breast
C1403582|T081|Observation of a mass
C1403582|T081|Molar Mass
C1403582|T081|Molecular Weights
C1403582|T081|Breast lump (finding)
C1403582|T081|Pulmonary Mass
C1403582|T081|MASS BREAST (NOS)
C1403582|T081|Superficial mass
C1403582|T081|Hepatic Mass
C1403582|T081|LIVER MASS
C1403582|T081|Liver mass
C1403582|T081|mass in or on skin
C1403582|T081|Liver Mass
C1403582|T081|breast mass
C1403582|T081|Superficial mass (finding)
C1403582|T081|Mass of body structure
C1403582|T081|Weight, Molecular
C1403582|T081|BREAST LUMPS
C1403582|T081|Molecular Mass
C1403582|T081|breast nodule
C1403582|T081|superficial mass
C1403582|T081|Lump in Breast
C1403582|T081|Lumpy breasts
C1403582|T081|Lump
C1403582|T081|density
C1403582|T081|Breast lump NOS
C1403582|T081|lung mass
C1403582|T081|LUNG MASS
C1403582|T081|breast density
C1403582|T081|Breast irregular nodularity
C1403582|T081|Breast nodule
C1403582|T081|BREAST NODULE
C1403582|T081|Mammary gland mass
C1403582|T081|molecular mass
C1403582|T081|Liver mass (finding)
C1403582|T081|nodular enhancement
C1403582|T081|extramammary mass
C1403582|T081|Localised mass
C1403582|T081|Breast lump
C1403582|T081|MW
C1709576|T033|Pleural Mass
C1511303|T191|Breast Carcinoma with Melanotic Features
CL412339|T061|Whole Breast Irradiation
CL412339|T061|whole breast irradiation
C0280401|T191|Recurrent Laryngeal Squamous Cell Carcinoma
C0280401|T191|Relapsed Larynx Squamous Cell Carcinoma
C0280401|T191|Relapsed Larynx Epidermoid Carcinoma
C0280401|T191|Recurrent Larynx Squamous Cell Carcinoma
C0280401|T191|Recurrent Larynx Epidermoid Carcinoma
C0280401|T191|Laryngeal squamous cell carcinoma recurrent
C0280401|T191|Relapsed Laryngeal Epidermoid Carcinoma
C0280401|T191|Recurrent Epidermoid Carcinoma of Larynx
C0280401|T191|Recurrent Squamous Cell Carcinoma of Larynx
C0280401|T191|Recurrent Laryngeal Epidermoid Carcinoma
C0280401|T191|Relapsed Squamous Cell Carcinoma of Larynx
C0280401|T191|epidermoid carcinoma of the larynx, recurrent
C0280401|T191|Relapsed Epidermoid Carcinoma of the Larynx
C0280401|T191|squamous cell carcinoma of the larynx, recurrent
C0280401|T191|Recurrent Epidermoid Carcinoma of the Larynx
C0280401|T191|Relapsed Laryngeal Squamous Cell Carcinoma
C0280401|T191|recurrent squamous cell carcinoma of the larynx
C0280401|T191|laryngeal squamous cell carcinoma, recurrent
C0280401|T191|Recurrent Squamous Cell Carcinoma of the Larynx
C0280401|T191|larynx squamous cell carcinoma, recurrent
C0280401|T191|Relapsed Epidermoid Carcinoma of Larynx
C0280401|T191|Relapsed Squamous Cell Carcinoma of the Larynx
C1831786|T061|Hypofractionated Radiation Therapy
C1831786|T061|hypofractionation
C1831786|T061|Hypofractionated Radiotherapy
C1831786|T061|hypofractionated radiation therapy
C1332623|T191|Breast Carcinoma Metastatic to the Bone
C0021308|T046|Ischemic Necrosis
C0021308|T046|avascular necrosis
C0021308|T046|Infarct (morphologic abnormality)
C0021308|T046|Ischemic necrosis
C0021308|T046|AVASCULAR NECROSIS
C0021308|T046|Avascular necrosis
C0021308|T046|Infarct
C0021308|T046|Infarction [Disease/Finding]
C0021308|T046|Avascular necrosis (morphologic abnormality)
C0021308|T046|NECROSIS ISCHEMIC
C0021308|T046|Infarcts
C0021308|T046|INFARCT
C0021308|T046|Necrosis, Avascular, of Bone
C0021308|T046|infarct
C0021308|T046|AVN - Avascular necrosis of bone
C0021308|T046|Bone Avascular Necrosis
C0021308|T046|ischemic necrosis
C0021308|T046|Avascular necrosis of bone
C0021308|T046|NECROSIS ISCHAEMIC
C0021308|T046|Infarction
C0021308|T046|Necrosis ischaemic
C0021308|T046|infarction
C0021308|T046|INFARCT INFARCTION
C0021308|T046|Avascular Necrosis of Bone
C0021308|T046|Ischaemic necrosis
C0021308|T046|Necrosis ischemic
C0021308|T046|Avascular Necrosis
C0021308|T046|avascular necrosis of bone
C0021308|T046|Avascular necrosis of bone (disorder)
C0021308|T046|Infarctions
C0021308|T046|Infarction NOS
C1332187|T191|Adult Brain Glioblastoma
C1332187|T191|Adult Brain Glioblastoma Multiforme
C0855010|T191|Recurrent Peripheral Primitive Neuroectodermal Tumor of Bone
C0855010|T191|Recurrent Neuroepithelioma of Bone
C0855010|T191|Recurrent PNET of Bone
C0424862|T033|Circumference of lump
C0424862|T033|Circumference of lump (observable entity)
C1334627|T191|TSH-Producing Pituitary Gland Carcinoma
C1334627|T191|Thyrotropin Producing Pituitary Gland Carcinoma
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Tumor of Pituitary Gland
C1334627|T191|Malignant TSH Producing Neoplasm of Pituitary Gland
C1334627|T191|Malignant TSH Producing Tumor of the Pituitary
C1334627|T191|Malignant TSH Secreting Neoplasm of Pituitary
C1334627|T191|Malignant Thyrotropinoma of Pituitary
C1334627|T191|Malignant Thyrotropinoma of the Pituitary
C1334627|T191|Malignant TSH Producing Pituitary Neoplasm
C1334627|T191|Malignant TSH Secreting Tumor of Pituitary Gland
C1334627|T191|Malignant TSH Producing Neoplasm of Pituitary
C1334627|T191|Malignant TSH Producing Pituitary Gland Tumor
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Neoplasm of the Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Tumor of the Pituitary
C1334627|T191|Malignant Thyrotropinoma of the Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Neoplasm of the Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Tumor
C1334627|T191|TSH Producing Pituitary Gland Carcinoma
C1334627|T191|Malignant Pituitary Gland Thyrotropinoma
C1334627|T191|Malignant TSH Producing Tumor of Pituitary Gland
C1334627|T191|Malignant TSH Producing Neoplasm of the Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Tumor of Pituitary
C1334627|T191|Malignant TSH Producing Pituitary Gland Neoplasm
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Pituitary Gland Tumor
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Tumor of Pituitary
C1334627|T191|Malignant TSH Producing Pituitary Tumor
C1334627|T191|Malignant TSH Secreting Pituitary Tumor
C1334627|T191|Malignant TSH Producing Neoplasm of the Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Tumor of the Pituitary Gland
C1334627|T191|Malignant TSH Producing Tumor of the Pituitary Gland
C1334627|T191|Malignant TSH Secreting Pituitary Gland Neoplasm
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Tumor of the Pituitary Gland
C1334627|T191|Malignant TSH Secreting Tumor of the Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Pituitary Gland Tumor
C1334627|T191|Malignant Pituitary Thyrotropinoma
C1334627|T191|Malignant TSH Producing Tumor of Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Pituitary Neoplasm
C1334627|T191|Malignant TSH Secreting Neoplasm of the Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Neoplasm of Pituitary
C1334627|T191|Malignant Thyrotropinoma
C1334627|T191|Malignant TSH Secreting Neoplasm of Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Pituitary Neoplasm
C1334627|T191|Malignant TSH Secreting Tumor of Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Pituitary Gland Neoplasm
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Neoplasm of Pituitary
C1334627|T191|Malignant TSH Secreting Tumor of the Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Neoplasm of the Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Neoplasm of the Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Tumor of Pituitary Gland
C1334627|T191|Malignant TSH Secreting Pituitary Neoplasm
C1334627|T191|Malignant Thyrotropinoma of Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Neoplasm of Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Neoplasm of Pituitary Gland
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Pituitary Gland Neoplasm
C1334627|T191|Malignant Thyroid Stimulating Hormone Producing Pituitary Tumor
C1334627|T191|Malignant TSH Secreting Neoplasm of the Pituitary Gland
C1334627|T191|Malignant TSH Secreting Pituitary Gland Tumor
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Tumor of the Pituitary
C1334627|T191|Malignant Thyroid Stimulating Hormone Secreting Pituitary Tumor
C1708069|T047|Flap Tissue Necrosis
C1708069|T047|NECROSIS OF FLAP TISSUE
C1708069|T047|FLAP TISSUE, NECROSIS OF
C1708069|T047|TISSUE, NECROSIS OF FLAP
C0475391|T185|T3b Stage Finding
C0475391|T185|T3b tumor stage
C0475391|T185|T3b
C0475391|T185|T3b Primary Tumor Finding
C0475391|T185|T3b Tumor Finding
C0475391|T185|T3b Cancer Stage Finding
C0475391|T185|T3b Primary Tumor Stage Finding
C0475391|T185|Tumor stage T3b
C0475391|T185|T3b TNM Finding
C0475391|T185|T3b Tumor Stage
C0475391|T185|Tumor Stage T3b
C0475391|T185|T3b Stage
C0475391|T185|Tumour stage T3b
C0475391|T185|Tumor stage T3b (finding)
C2825182|T061|Atrial Ablation
C2825182|T061|ABLATION, ATRIAL
C1335258|T191|PRETEXT Stage 4 Hepatoblastoma
C2732473|T191|Microinvasive Breast Carcinoma
C2732473|T191|Ductal Carcinoma In Situ with Microinvasion
C2732473|T191|MIC
C2732473|T191|Ductal carcinoma in situ with microinvasion (morphologic abnormality)
C2732473|T191|DCISM
C2732473|T191|Ductal carcinoma in situ with microinvasion
C1335714|T191|Recurrent Metastatic Squamous Cell Carcinoma to the Neck with Occult Primary
C1335714|T191|Relapsed Metastatic Squamous Cell Carcinoma to the Neck with Occult Primary
C1335714|T191|Relapsed Metastatic Epidermoid Carcinoma to the Neck with Occult Primary
C1335714|T191|Relapsed Metastatic Squamous Cell Neck Cancer with Occult Primary
C1335714|T191|Recurrent Metastatic Squamous Cell Cancer to the Neck with Occult Primary
C1335714|T191|Recurrent Metastatic Epidermoid Carcinoma to the Neck with Occult Primary
C0854802|T191|Recurrent Chronic Lymphocytic Leukemia
C0854802|T191|leukemia, relapsed chronic lymphocytic
C0854802|T191|Relapsed Chronic Lymphoid Leukemia
C0854802|T191|Chronic lymphocytic leukaemia recurrent
C0854802|T191|chronic lymphocytic leukemia, relapsed
C0854802|T191|Recurrent Chronic Lymphoid Leukemia
C0854802|T191|Relapsed Chronic Lymphocytic Leukemia
C0854802|T191|relapsed CLL
C0854802|T191|Recurrent Chronic Lymphogenous Leukemia
C0854802|T191|CLL, relapsed
C0854802|T191|Chr lymp leuk in relapse
C0854802|T191|Chronic lymphocytic leukemia recurrent
C0854802|T191|relapsed chronic lymphocytic leukemia
C0854802|T191|Chronic lymphoid leukemia, in relapse
C0854802|T191|lymphocytic leukemia, relapsed chronic
C0854802|T191|Relapsed Chronic Lymphogenous Leukemia
C0854802|T191|Chronic Lymphocytic Leukemia Recurrent
C1334731|T191|Metastatic Malignant Neoplasm to the Nasopharynx
C1334731|T191|Metastatic Tumor to the Nasopharynx
C1334731|T191|Metastasis to the Nasopharynx
C1334731|T191|Metastatic Neoplasm to the Nasopharynx
C0854989|T191|Recurrent Squamous Cell Lung Carcinoma
C0854989|T191|Recurrent Squamous Cell Carcinoma of the Lung
C0854989|T191|Recurrent Squamous Cell Carcinoma of Lung
C0854989|T191|Lung squamous cell carcinoma recurrent
C0280191|T191|Recurrent Adult Lymphoblastic Lymphoma
C0280191|T191|Recurrent Adult Precursor Lymphoblastic Lymphoma
C0280191|T191|recurrent adult lymphoblastic lymphoma
C0280191|T191|adult lymphoblastic lymphoma, relapsed
C0280191|T191|lymphoblastic lymphoma, adult, recurrent
C0280191|T191|Adult Recurrent Lymphoblastic Lymphoma
C0280191|T191|relapsed adult lymphoblastic lymphoma
C0280191|T191|lymphoblastic lymphoma, recurrent, adult
C0280191|T191|adult lymphoblastic lymphoma, recurrent
C0279766|T034|Progesterone Receptor Negative
C0279766|T034|PR-
C0279766|T034|negative progesterone receptor
C0279766|T034|progesterone receptor negative
C2986680|T191|Stage IV Childhood Non-Hodgkin Lymphoma
C2986680|T191|stage IV childhood non-Hodgkin lymphoma
C0144576|T121|Paclitaxel
C0144576|T121|PACLITAXEL
C0144576|T121|5Beta,20-epoxy-1,2alpha,4,7beta,10beta,13alpha-hexahydroxytax-11-en-9-one, 4,10-Diacetate 2-Benzoate 13-Ester with (2R,3S)-N-Benzoyl-3-phenylisoserine
C0144576|T121|Taxol
C0144576|T121|Bristaxol
C0144576|T121|Taxol Konzentrat
C0144576|T121|Anzatax
C0144576|T121|Asotax
C0144576|T121|[2aR-[2a Alpha,4beta,4a beta,6beta,9alpha(alphaR*,betaS*),-11alpha,12alpha,12a alpha,12b alpha]]-beta-(benzoylamino)-alpha-hydroxybenzene-propanoic acid 6,12b-bis(acetyloxy)-12-(benzoyloxy)-1a,33,4,-41,5,6,9,10,11,12,12a,12b-dodecahydro-4,11-dihydroxy-41,8,-12,13-tetramethyl-5-oxo-7,11-methano-1H-cyclodeca[3,4]benz[1,2-b]oxet-9-yl Ester
C0144576|T121|Praxel
C0144576|T121|paclitaxel
CL376186|T191|Recurrent Childhood Non-Hodgkin Lymphoma
C1321211|T033|Tumor nodule size, additional dimension
C1321211|T033|Tumor nodule size, additional dimension (observable entity)
C1321211|T033|Tumour nodule size, additional dimension
C1334797|T191|Monomorphic B-Cell Post-Transplant Lymphoproliferative Disorder
C1334797|T191|Monomorphic B-Cell PTLD
C0863127|T191|Chemotherapy-Related Leukemia
C0863127|T191|Leukemia secondary to oncology chemotherapy
CL388374|T061|Accelerated Partial Breast Irradiation
CL388374|T061|APBI
CL388374|T061|accelerated partial breast irradiation
C1333381|T033|Encapsulated Mass
C1333381|T033|Encapsulated
C1333381|T033|encapsulated
C1300500|T201|Tumor size, dominant nodule, additional dimension, in specimen obtained by prostatic enucleation
C1300500|T201|Tumour size, dominant nodule, additional dimension, in specimen obtained by prostatic enucleation
C1300500|T201|Tumor size, dominant nodule, additional dimension, in specimen obtained by prostatic enucleation (observable entity)
C1336863|T191|Undifferentiated Prostate Carcinoma
C1336863|T191|Undifferentiated Prostatic Carcinoma
C1336863|T191|Undifferentiated Carcinoma of the Prostate
C1336863|T191|Undifferentiated Carcinoma of Prostate
C0877578|T191|Therapy-Related Malignant Neoplasm
C0877578|T191|Therapy Related Cancer
C0877578|T191|Therapy Related Malignant Neoplasm
C0877578|T191|Treatment related secondary malignancy
C0877578|T191|Iatrogenic Cancer
C0877578|T191|Therapy Related Malignant Tumor
C1336769|T191|Topoisomerase II Inhibitor-Related Acute Myeloid Leukemia
C1336769|T191|Topoisomerase II Inhibitor-Related AML
C1336769|T191|Topoisomerase II Inhibitor Related Acute Myeloid Leukemia
C1273121|T081|Polyp stalk length
C1273121|T081|Polyp stalk length (observable entity)
C0334384|T191|Invasive Ductal and Lobular Carcinoma In Situ
C0334384|T191|Lobular Carcinoma in situ and Infiltrating Ductal Carcinoma
C0334384|T191|Lobular Carcinoma in situ and Invasive Ductal Carcinoma
C0334384|T191|LCIS and Infiltrating Ductal Carcinoma
C0334384|T191|Infiltrating Ductal and Lobular Carcinoma in situ
C1708790|T033|Lymphatic Invasion
C1708790|T033|Lymphovascular Invasion
C0445037|T033|M1c Stage Finding
C0445037|T033|Metastasis stage M1c (finding)
C0445037|T033|M1c Cancer Stage Finding
C0445037|T033|M1c Distant Metastasis Stage Finding
C0445037|T033|M1c Metastasis Finding
C0445037|T033|M1c Stage
C0445037|T033|Metastasis Stage M1c
C0445037|T033|M1c TNM Finding
C0445037|T033|M1c Metastasis Stage
C0445037|T033|Metastasis stage M1c
C0445037|T033|M1c
C0445037|T033|M1c Distant Metastasis Finding
C1334285|T191|Ionizing Radiation-Related Malignant Neoplasm
C1708784|T191|Lung Spindle Cell Carcinoma
CL433931|T061|Percutaneous Cryosurgery
CL433931|T061|percutaneous cryosurgery
C0334271|T191|Sarcomatoid Transitional Cell Carcinoma
C0334271|T191|Transitional cell carcinoma, spindle cell
C0334271|T191|Transitional cell carcinoma - spindle cell
C0334271|T191|Transitional Spindle Cell Carcinoma
C0334271|T191|Transitional cell carcinoma, spindle cell (morphologic abnormality)
C0334271|T191|Transitional cell carcinoma, sarcomatoid
C0334271|T191|Transitional Cell Spindle Cell Carcinoma
CL433972|T191|Familial Neuroblastoma
CL433972|T191|Hereditary Neuroblastoma
CL433972|T191|hereditary neuroblastoma
CL433972|T191|neuroblastoma, hereditary
C0475371|T033|T0 stage
C0475371|T033|T0 Cancer Stage Finding
C0475371|T033|T0
C0475371|T033|T0 Tumor Finding
C0475371|T033|T0 Stage Finding
C0475371|T033|T0 Stage
C0475371|T033|Tumor Stage T0
C0475371|T033|T0 category (finding)
C0475371|T033|T0 category
C0475371|T033|T0 Primary Tumor Finding
C0475371|T033|T0 Tumor Stage
C0475371|T033|Tumour stage T0
C0475371|T033|T0 TNM Finding
C0475371|T033|T0 Primary Tumor Stage Finding
C0475371|T033|Tumor stage T0
CL414453|T191|Childhood Anaplastic Astrocytoma
CL414453|T191|Grade III Pediatric Astrocytic Neoplasm
CL414453|T191|astrocytoma, grade III childhood
CL414453|T191|grade III pediatric astrocytic tumor
CL414453|T191|undifferentiated pediatric astrocytoma
CL414453|T191|Undifferentiated Childhood Astrocytoma
CL414453|T191|grade III childhood astrocytic neoplasm
CL414453|T191|pediatric anaplastic astrocytoma
CL414453|T191|undifferentiated childhood astrocytoma
CL414453|T191|Grade III Childhood Astrocytic Tumor
CL414453|T191|Anaplastic Childhood Astrocytoma
CL414453|T191|grade III childhood astrocytic tumor
CL414453|T191|Grade III Pediatric Astrocytoma
CL414453|T191|Grade III Childhood Astrocytoma
CL414453|T191|anaplastic astrocytoma, childhood
CL414453|T191|anaplastic childhood astrocytoma
CL414453|T191|Undifferentiated Pediatric Astrocytoma
CL414453|T191|Grade III Childhood Astrocytic Neoplasm
CL414453|T191|Grade III Pediatric Astrocytic Tumor
CL414453|T191|Anaplastic Pediatric Astrocytoma
CL414453|T191|grade III pediatric astrocytoma
CL414453|T191|grade III pediatric astrocytic neoplasm
CL414453|T191|anaplastic pediatric astrocytoma
CL414453|T191|childhood anaplastic astrocytoma
CL414453|T191|astrocytoma, childhood anaplastic
CL414453|T191|grade III childhood astrocytoma
C1334276|T191|Invasive Ductal and Invasive Lobular Breast Carcinoma
C1334276|T191|Infiltrating Ductal and Infiltrating Lobular Breast Carcinoma
C1332988|T191|Childhood Ovarian Dysgerminoma
C1332988|T191|Pediatric Ovarian Dysgerminoma
C0855002|T191|Recurrent Lung Carcinoma
C0855002|T191|Lung cancer recurrent
C0855002|T191|Relapsed Unspecified Lung Carcinoma
C0855002|T191|Recurrent Unspecified Lung Carcinoma
C0855002|T191|Relapsed Unspecified Carcinoma of Lung
C0855002|T191|Pulmonary carcinoma recurrent
C0855002|T191|Lung carcinoma cell type unspecified recurrent
C0855002|T191|Pulmonary carcinoma cell type unspecified recurrent
C0855002|T191|Recurrent Lung Cancer
C0855002|T191|Relapsed Unspecified Carcinoma of the Lung
C0855002|T191|Cancer of lung recurrent
C0855002|T191|Lung carcinoma recurrent
C0855002|T191|Recurrent Unspecified Carcinoma of Lung
C0855002|T191|Recurrent Unspecified Carcinoma of the Lung
C0475397|T185|T4c Stage Finding
C0475397|T185|T4c Stage
C0475397|T185|Tumor stage T4c
C0475397|T185|T4c
C0475397|T185|T4c Tumor Finding
C0475397|T185|T4c Cancer Stage Finding
C0475397|T185|T4c Primary Tumor Stage Finding
C0475397|T185|T4c TNM Finding
C0475397|T185|Tumour stage T4c
C0475397|T185|T4c Tumor Stage
C0475397|T185|Tumor Stage T4c
C0475397|T185|T4c Primary Tumor Finding
C0475397|T185|Tumor stage T4c (finding)
C1292776|T191|Therapy-Related Myeloid Neoplasm
C1292776|T191|Therapy-Related AML and MDS
C1292776|T191|Therapy-Related Acute Myeloid Leukemia and Myelodysplastic Syndrome
C1292776|T191|Acute Myeloid Leukaemias and Myelodysplastic Syndromes, Therapy-Related
C1335700|T191|Recurrent Female Reproductive System Carcinoma
C1335700|T191|Recurrent Female Reproductive System Cancer
C1333085|T191|Colon Carcinoma Metastatic to the Liver
C1332638|T191|Breast Small Cell Carcinoma
C1332638|T191|Oat Cell Carcinoma of Breast
C1332638|T191|Mammary Small Cell Carcinoma
C1332638|T191|Small Cell Carcinoma of the Breast
C1332638|T191|Small Cell Neuroendocrine Carcinoma of the Breast
C1332638|T191|Oat Cell Carcinoma of the Breast
C1332638|T191|Small Cell Neuroendocrine Carcinoma of Breast
C1332638|T191|Small Cell Carcinoma of Breast
C0457423|T033|V2 Cancer Stage Finding
C0457423|T033|V2
C0457423|T033|V2 stage
C0457423|T033|V2: macroscopic venous invasion
C0457423|T033|V2 Venous Stage
C0457423|T033|Venous stage V2
C0457423|T033|V2 Stage
C0457423|T033|Venous Stage V2
C0457423|T033|V2 Venous Invasion Finding
C0457423|T033|V2 Stage Finding
C0457423|T033|V2 TNM Finding
C0457423|T033|V2 stage (finding)
C115441|T191|Recurrent Primary Peritoneal Carcinoma
C0854820|T191|Recurrent Anaplastic Large Cell Lymphoma
C0854820|T191|Relapsed Anaplastic Large Cell Lymphoma
C0854820|T191|Anaplastic large cell lymphoma T- and null-cell types recurrent
C100079|T002|Tobacco Smoking
C100079|T002|Smoking Tobacco
C100079|T002|Smoke
C100079|T002|tobacco smoke
C100079|T002|Smoked Tobacco
C100079|T002|Tobacco Smoke
C100079|T002|Smoking
C100079|T002|Tobacco smoke
C100079|T002|Tobacco smoke (substance)
C0281605|T061|Bone Marrow Ablation with Stem Cell Support
C0449712|T082|Pituitary adenoma size
C0449712|T082|Pituitary adenoma size (observable entity)
C0449712|T082|Size of pituitary adenoma
C0279758|T034|Estrogen Receptor Status Unknown
C0279758|T034|estrogen receptor status unknown
C0279758|T034|Unknown Status, Estrogen Receptor
C0279758|T034|unknown status, estrogen receptor
C0855186|T191|Recurrent Bladder Squamous Cell Carcinoma
C0855186|T191|Squamous cell bladder carcinoma recurrent
C0855186|T191|Relapsed Squamous Cell Carcinoma of the Urinary Bladder
C0855186|T191|Relapsed Urinary Bladder Squamous Cell Carcinoma
C0855186|T191|Relapsed Squamous Cell Carcinoma of the Bladder
C0855186|T191|Squamous cell carcinoma of the bladder recurrent
C0855186|T191|Recurrent Urinary Bladder Epidermoid Carcinoma
C0855186|T191|Squamous Cell Carcinoma of the Bladder, Recurrent
C0855186|T191|Relapsed Bladder Epidermoid Carcinoma
C0855186|T191|Relapsed Epidermoid Carcinoma of the Bladder
C0855186|T191|Bladder squamous cell carcinoma recurrent
C0855186|T191|Relapsed Bladder Squamous Cell Carcinoma
C0855186|T191|Relapsed Epidermoid Carcinoma of Urinary Bladder
C0855186|T191|Recurrent Epidermoid Carcinoma of the Bladder
C0855186|T191|Relapsed Epidermoid Carcinoma of Bladder
C0855186|T191|Recurrent Epidermoid Carcinoma of Urinary Bladder
C0855186|T191|Squamous Cell Carcinoma of Bladder, Recurrent
C0855186|T191|Recurrent Squamous Cell Carcinoma of Bladder
C0855186|T191|Relapsed Epidermoid Carcinoma of the Urinary Bladder
C0855186|T191|Relapsed Squamous Cell Carcinoma of Bladder
C0855186|T191|Recurrent Squamous Cell Carcinoma of the Urinary Bladder
C0855186|T191|Recurrent Epidermoid Carcinoma of Bladder
C0855186|T191|Relapsed Urinary Bladder Epidermoid Carcinoma
C0855186|T191|Recurrent Squamous Cell Carcinoma of the Bladder
C0855186|T191|Recurrent Epidermoid Carcinoma of the Urinary Bladder
C0855186|T191|Relapsed Squamous Cell Carcinoma of Urinary Bladder
C0855186|T191|Recurrent Urinary Bladder Squamous Cell Carcinoma
C0855186|T191|Recurrent Bladder Epidermoid Carcinoma
C0855186|T191|Recurrent Squamous Cell Carcinoma of Urinary Bladder
C1705427|T049|Germline Mutation Abnormality
C1705427|T049|Germline Mutation
C115442|T191|Recurrent Lip and Oral Cavity Squamous Cell Carcinoma
C1272779|T201|Tumor size, largest dimension
C1272779|T201|Tumor size, greatest dimension
C1272779|T201|Tumor size, largest dimension (observable entity)
C1272779|T201|Tumour size, greatest dimension
C1272779|T201|Tumour size, largest dimension
C3272818|T191|Colorectal Sarcomatoid Carcinoma
C3272818|T191|Colorectal Spindle Cell Carcinoma
C1332999|T191|Childhood Primary Cutaneous Anaplastic Large Cell Lymphoma
C1332999|T191|Pediatric Primary Cutaneous K-1+ Anaplastic Large Cell Lymphoma
C1332999|T191|Childhood Primary Cutaneous CD30-Positive Anaplastic Large Cell Lymphoma
C1332999|T191|Childhood Primary Cutaneous CD30+ Anaplastic Large Cell Lymphoma
C1332999|T191|Childhood Primary Cutaneous Ki-1+ Anaplastic Large Cell Lymphoma
C1332999|T191|Childhood Primary Cutaneous Ki-1 Positive Anaplastic Large Cell Lymphoma
C1332999|T191|Pediatric Primary Cutaneous CD30+ Anaplastic Large Cell Lymphoma
C1332999|T191|Pediatric Primary Cutaneous Anaplastic Large Cell Lymphoma
C0854796|T191|Non-Resectable Hepatoblastoma
C0854796|T191|Hepatoblastoma, Nonresectable
C0854796|T191|Unresectable Hepatoblastoma
C1709108|T033|N3a Stage Finding
C1709108|T033|N3a Regional Lymph Node Stage Finding
C1709108|T033|N3a Node Finding
C1709108|T033|N3a Cancer Stage Finding
C1709108|T033|N3a Stage
C1709108|T033|N3a TNM Finding
C1709108|T033|N3a
C1709108|T033|N3a Node Stage
C1709108|T033|N3a Lymph Node Finding
C1709108|T033|Lymph Node Stage N3a
C1709108|T033|N3a Regional Lymph Nodes Finding
C1709108|T033|Node Stage N3a
C1709108|T033|N3a Lymph Node Stage
C0862642|T191|Stage III Prostate Adenocarcinoma
C0862642|T191|Stage III Prostate Adenocarcinoma AJCC v7
C1334822|T033|Multinodular Mass
C1333179|T191|Cutaneous Radiation-Related Angiosarcoma
C1333179|T191|Cutaneous Radiation-Induced Angiosarcoma
C0280733|T191|Recurrent Carcinoma of Unknown Primary
C1512032|T049|Dominant-Negative Mutation
C1512032|T049|Dominant-Negative Mutant
C1512032|T049|Dominant-Negative Mutation Abnormality
C1512032|T049|Dominant Negative
CL343570|T191|Childhood Supratentorial Primitive Neuroectodermal Tumor
CL343570|T191|supratentorial primitive neuroectodermal tumor, childhood
CL343570|T191|Brain tumor, child: PNET
CL343570|T191|childhood supratentorial PNET
CL343570|T191|PNET, supratentorial, pediatric
CL343570|T191|childhood supratentorial primitive neuroectodermal tumor
CL343570|T191|PNET, pediatric supratentorial
CL343570|T191|neuroectodermal tumor, pediatric, primitive, supratentorial
CL343570|T191|primitive neuroectodermal tumor, supratentorial, pediatric
CL343570|T191|pediatric supratentorial primitive neuroectodermal tumor
CL343570|T191|primitive neuroectodermal tumor, childhood supratentorial
CL343570|T191|pediatric primitive neuroectodermal tumor, supratentorial
CL343570|T191|supratentorial primitive neuroectodermal tumor, pediatric
CL343570|T191|pediatric supratentorial PNET
CL343570|T191|PNET, supratentorial, childhood
CL343570|T191|PNET, childhood supratentorial
CL343570|T191|primitive neuroectodermal tumor, pediatric supratentorial
CL343570|T191|neuroectodermal tumor, childhood, primitive, supratentorial
CL343570|T191|childhood primitive neuroectodermal tumor, supratentorial
CL343570|T191|primitive neuroectodermal tumor, supratentorial, childhood
C1332279|T191|Anaplastic Brain Stem Astrocytoma
C1332279|T191|Anaplastic Brainstem Astrocytoma
CL376163|T191|Recurrent Extragonadal Seminoma
CL376163|T191|recurrent extragonadal seminoma
C1708349|T191|Hereditary Diffuse Gastric Adenocarcinoma
C1708349|T191|gastric cancer, hereditary diffuse
C1708349|T191|gastric cancer, familial
C1708349|T191|HDGC
C1708349|T191|hereditary diffuse gastric cancer
C1708349|T191|GASTRIC CANCER, FAMILIAL DIFFUSE
C1708349|T191|familial gastric cancer
C1708349|T191|GASTRIC CANCER, HEREDITARY DIFFUSE
C1708349|T191|Hereditary Diffuse Gastric Cancer
C1708349|T191|Gastric Cancer, Familial Diffuse
C1512744|T191|Infiltrating Bladder Urothelial Carcinoma, Sarcomatoid Variant with Heterologous Elements
C1514588|T033|Pseudopalisading Necrosis
C1332993|T191|Childhood Ovarian Yolk Sac Tumor
C1332993|T191|Pediatric Ovarian Yolk Sac Tumor
C1332993|T191|Childhood Ovarian Endodermal Sinus Tumor
C1332993|T191|Childhood Ovarian Yolk Sac Neoplasm
C1332993|T191|Pediatric Ovarian Endodermal Sinus Tumor
C1332993|T191|Pediatric Ovarian Endodermal Sinus Neoplasm
C1332993|T191|Childhood Ovarian Endodermal Sinus Neoplasm
C1332993|T191|Pediatric Ovarian Yolk Sac Neoplasm
C1300513|T201|Tumor size, invasive component
C1300513|T201|Tumor size, invasive component (observable entity)
C1300513|T201|Tumour size, invasive component
C1336810|T191|Transplant-Related Hematologic Malignancy
C1512748|T191|Infiltrating Bladder Urothelial Carcinoma with Squamous Differentiation
C1512748|T191|Infiltrating Bladder Urothelial Carcinoma with Squamous
C1332610|T191|Brain Stem Glioblastoma
C1332610|T191|Glioblastoma Multiforme of Brainstem
C1332610|T191|Grade IV Brainstem Astrocytic Neoplasm
C1332610|T191|Grade IV Astrocytic Neoplasm of the Brainstem
C1332610|T191|Grade IV Brain Stem Astrocytic Tumor
C1332610|T191|Glioblastoma Multiforme of the Brain Stem
C1332610|T191|Grade IV Brain Stem Astrocytic Neoplasm
C1332610|T191|Glioblastoma Multiforme of Brain Stem
C1332610|T191|Brain Stem Glioblastoma Multiforme
C1332610|T191|Grade IV Astrocytic Tumor of the Brain Stem
C1332610|T191|Grade IV Astrocytic Tumor of Brain Stem
C1332610|T191|Grade IV Astrocytic Tumor of the Brainstem
C1332610|T191|Grade IV Astrocytic Neoplasm of Brain Stem
C1332610|T191|Grade IV Astrocytic Tumor of Brainstem
C1332610|T191|Brainstem Glioblastoma
C1332610|T191|Grade IV Astrocytic Neoplasm of Brainstem
C1332610|T191|Glioblastoma Multiforme of the Brainstem
C1332610|T191|Grade IV Astrocytic Neoplasm of the Brain Stem
C1332610|T191|Grade IV Brainstem Astrocytic Tumor
C1332610|T191|Brainstem Glioblastoma Multiforme
C1519560|T201|Total Nodal Irradiation
C1519560|T201|total nodal irradiation
C1519560|T201|total lymphoid irradiation
C1519560|T201|TLI
C0278321|T061|Bilateral Oophorectomy
C0278321|T061|Female Castration
C0278321|T061|Ovariectomies, Bilateral
C0278321|T061|Female Castrations
C0278321|T061|Oophorectomy bilateral
C0278321|T061|Oth remove both ovaries
C0278321|T061|Other removal of both ovaries at same operative episode
C0278321|T061|Castration, Female
C0278321|T061|Bilateral oophorectomy (procedure)
C0278321|T061|Bilateral Ovariectomy
C0278321|T061|Castrations, Female
C0278321|T061|Ovariectomy, Bilateral
C0278321|T061|Spay operation
C0278321|T061|Bilateral oophorectomy
C0278321|T061|Female castration
C0278321|T061|Bilateral Ovariectomies
C1705057|T201|Circumferential Resection Margin
C1705057|T201|CRM
C2827060|T033|Polyp Tip
C0220612|T191|Childhood Non-Hodgkin Lymphoma
C0220612|T191|Pediatric Non-Hodgkin Lymphoma
C0220612|T191|Childhood Non-Hodgkin's Lymphoma
C0220612|T191|Pediatric Non-Hodgkin's Lymphoma
C0279083|T191|Meningeal Chronic Myelogenous Leukemia, BCR-ABL1 Positive
C0279083|T191|Meningeal Chronic Myelogenous Leukemia
C0855008|T191|Metastatic Peripheral Primitive Neuroectodermal Tumor of Bone
C0855008|T191|Metastatic Peripheral Neuroepithelioma of Bone
C1332079|T191|Anaplastic Large Cell Lymphoma, ALK-Positive
C1332079|T191|ALKoma
C1332079|T191|ALCL, ALK+
C1332079|T191|ALK-Positive Anaplastic Large Cell Lymphoma
C0279614|T191|Childhood Anaplastic Rhabdomyosarcoma
C0279614|T191|rhabdomyosarcoma, pediatric pleomorphic
C0279614|T191|rhabdomyosarcoma, childhood pleomorphic
C0279614|T191|childhood rhabdomyosarcoma, pleomorphic
C0279614|T191|Pleomorphic Childhood Rhabdomyosarcoma
C0279614|T191|pediatric rhabdomyosarcoma, pleomorphic
C0279614|T191|rhabdomyosarcoma, pleomorphic childhood
C0279614|T191|pleomorphic childhood rhabdomyosarcoma
C0279614|T191|Childhood Pleomorphic Rhabdomyosarcoma
C0279614|T191|Pediatric Pleomorphic Rhabdomyosarcoma
C0279614|T191|pleomorphic pediatric rhabdomyosarcoma
C1947968|T191|Carcinoma Metastatic to the Skin
C1947968|T191|Metastatic Skin Cancer
C1947968|T191|Metastatic Skin Carcinoma
C1335444|T191|Poorly Differentiated Malignant Neoplasm
C1706790|T191|Ameloblastic Carcinoma-Secondary Type (Dedifferentiated), Peripheral
C1706790|T191|Peripheral Ameloblastic Carcinoma
C0475383|T185|Tumor stage T1a
C0475383|T185|Tumor Stage T1a
C0475383|T185|T1a Stage
C0475383|T185|Tumor stage T1a (finding)
C0475383|T185|T1a Cancer Stage Finding
C0475383|T185|Tumour stage T1a
C0475383|T185|T1a Tumor Finding
C0475383|T185|T1a Primary Tumor Finding
C0475383|T185|T1a Stage Finding
C0475383|T185|T1a Primary Tumor Stage Finding
C0475383|T185|T1a
C0475383|T185|T1a TNM Finding
C0475383|T185|T1a Tumor Stage
C0441474|T061|Chemical Ablation
C0441474|T061|Chemical ablation
C0441474|T061|Chemical destruction
C0441474|T061|Chemical destruction (qualifier value)
C0441474|T061|ABLATION, CHEMICAL
C0950521|T061|CMF Regimen
C0950521|T061|CMF regimen
C0950521|T061|CMF
C0950521|T061|CTX/5-FU/MTX
C0950521|T061|Cytoxan-Methotrexate-Fluorouracil Regimen
C0950521|T061|Cyclophosphamide/Fluorouracil/Methotrexate
C0950521|T061|Cyclophosphamide-Methotrexate-Fluorouracil regimen
C1333982|T191|Hepatoblastoma with Pure Fetal Epithelial Differentiation
C1272618|T033|Polyp size, largest dimension
C1272618|T033|Polyp size greatest dimension
C1272618|T033|Polyp size, greatest dimension
C1272618|T033|Polyp size, largest dimension (observable entity)
C1332946|T191|Childhood Botryoid-Type Embryonal Rhabdomyosarcoma of the Vulva
C1332946|T191|Vulvar Childhood Botryoid-Type Embryonal Rhabdomyosarcoma
C1332946|T191|Childhood Sarcoma Botryoides of the Vulva
C1335719|T191|Recurrent Peripheral Primitive Neuroectodermal Tumor
C0886483|T191|Childhood Malignant Ovarian Germ Cell Tumor
C0886483|T191|childhood malignant ovarian germ cell tumor
C0278838|T191|Recurrent Prostate Carcinoma
C0278838|T191|Recurrent Prostate Cancer
C0278838|T191|recurrent prostate cancer
C0278838|T191|prostate cancer, recurrent
C0278838|T191|Carcinoma of the prostate recurrent
C0278838|T191|Recurrent Cancer of the Prostate
C0278838|T191|Recurrent Cancer of Prostate
C0278838|T191|Prostatic cancer recurrent
C0278838|T191|Prostate cancer recurrent
C1514513|T191|Prostate Ductal Adenocarcinoma, Solid Pattern
C1880568|T061|Ethanol Ablation Therapy
C1880568|T061|ethanol ablation
C1880568|T061|PEI
C1880568|T061|percutaneous ethanol injection
C1880568|T061|ethanol ablation therapy
C1880568|T061|alcohol ablation
C0861556|T191|Recurrent Oral Cavity Squamous Cell Carcinoma
C0861556|T191|Relapsed Epidermoid Carcinoma of Mouth
C0861556|T191|Recurrent Squamous Cell Carcinoma of the Mouth
C0861556|T191|Squamous cell carcinoma of the oral cavity recurrent
C0861556|T191|Relapsed Mouth Squamous Cell Carcinoma
C0861556|T191|Recurrent Squamous Cell Carcinoma of the Oral Cavity
C0861556|T191|Recurrent Epidermoid Carcinoma of the Mouth
C0861556|T191|Recurrent Squamous Cell Carcinoma of Oral Cavity
C0861556|T191|Recurrent Mouth Epidermoid Carcinoma
C0861556|T191|Relapsed Squamous Cell Carcinoma of the Mouth
C0861556|T191|Relapsed Epidermoid Carcinoma of Oral Cavity
C0861556|T191|Relapsed Epidermoid Carcinoma of the Mouth
C0861556|T191|Relapsed Squamous Cell Carcinoma of Oral Cavity
C0861556|T191|Recurrent Oral Cavity Epidermoid Carcinoma
C0861556|T191|Relapsed Epidermoid Carcinoma of the Oral Cavity
C0861556|T191|Recurrent Epidermoid Carcinoma of the Oral Cavity
C0861556|T191|Relapsed Mouth Epidermoid Carcinoma
C0861556|T191|Recurrent Squamous Cell Carcinoma of Mouth
C0861556|T191|Recurrent Epidermoid Carcinoma of Oral Cavity
C0861556|T191|Relapsed Squamous Cell Carcinoma of Mouth
C0861556|T191|Relapsed Oral Cavity Epidermoid Carcinoma
C0861556|T191|Relapsed Squamous Cell Carcinoma of the Oral Cavity
C0861556|T191|Recurrent Mouth Squamous Cell Carcinoma
C0861556|T191|Relapsed Oral Cavity Squamous Cell Carcinoma
C0861556|T191|Recurrent Epidermoid Carcinoma of Mouth
C0178421|T191|Fibroadenoma
C0178421|T191|BREAST, ADENOFIBROMA
C0178421|T191|BREAST FIBROADENOMA
C0178421|T191|BREAST, FIBROADENOMA
C0178421|T191|Breast Fibroadenoma
C0178421|T191|Fibroadenoma, no ICD-O subtype (morphologic abnormality)
C0178421|T191|Fibroadenoma of breast (disorder)
C0178421|T191|Fibroadenoma of breast
C0178421|T191|Breast mouse
C0178421|T191|FIBROADENOMA OF THE BREAST
C0178421|T191|Fibroadenoma [Disease/Finding]
C0178421|T191|Fibroadenoma, no ICD-O subtype
C0178421|T191|Breast fibroadenomas
C0178421|T191|Fibroadenoma, NOS
C0178421|T191|fibroadenoma
C0178421|T191|fibroadenoma of breast
C0178421|T191|Fibroadenomas
C0178421|T191|Fibroadenoma of Breast
C0178421|T191|FIBROADENOMA OF BREAST
C0178421|T191|Fibroadenoma of the Breast
C0178421|T191|FIBROADENOMA, BENIGN
C0281342|T061|Bone Marrow Ablation
C0281342|T061|bone marrow ablation
C0029936|T061|Oophorectomy
C0029936|T061|Female Castration
C0029936|T061|Ovary removal
C0029936|T061|Oophorectomy (procedure)
C0029936|T061|Ovariectomies
C0029936|T061|female gonadectomy
C0029936|T061|ovariectomy
C0029936|T061|OOPHORECTOMY
C0029936|T061|Excision of ovary
C0029936|T061|Oophorectomies
C0029936|T061|Ovariectomy
C0029936|T061|female castration
C0029936|T061|oophorectomy
C0029936|T061|Oophorectomy NOS
C0346989|T191|Metastatic Malignant Neoplasm to the Peritoneum
C0346989|T191|Metastases to peritoneum, NOS
C0346989|T191|Metastatic Neoplasm to the Peritoneum
C0346989|T191|Metastasis to the Peritoneum
C0149736|T033|Neck Mass
C0149736|T033|Mass of neck (finding)
C0149736|T033|Lump on neck
C0149736|T033|Mass of neck
C0149736|T033|NECK MASS
C0149736|T033|Neck Lump
C0149736|T033|Neck mass
C0279975|T191|Recurrent Ovarian Germ Cell Tumor
C0279975|T191|recurrent ovarian germ cell tumor
C0279975|T191|Recurrent Germ Cell Tumor of Ovary
C0279975|T191|Recurrent Germ Cell Neoplasm of Ovary
C0279975|T191|Relapsed Germ Cell Tumor of the Ovary
C0279975|T191|Relapsed Germ Cell Tumor of Ovary
C0279975|T191|Relapsed Ovarian Germ Cell Tumor
C0279975|T191|Relapsed Germ Cell Neoplasm of Ovary
C0279975|T191|Recurrent Ovarian Germ Cell Neoplasm
C0279975|T191|germ cell tumor, ovarian, recurrent
C0279975|T191|Recurrent Germ Cell Tumor of the Ovary
C0279975|T191|ovarian germ cell tumor, recurrent
C0279975|T191|Relapsed Ovarian Germ Cell Neoplasm
C0279975|T191|Recurrent Germ Cell Neoplasm of the Ovary
C0279975|T191|Relapsed Germ Cell Neoplasm of the Ovary
C0854823|T191|Stage II Anaplastic Large Cell Lymphoma
C0854823|T191|Anaplastic Large Cell Lymphoma Stage II
C0854823|T191|Anaplastic Large Cell Lymphoma T- and Null-Cell Types Stage II
C3273216|T191|Invasive Lobular Breast Carcinoma, Pleomorphic Variant
C2985392|T061|Argon Beam Coagulator Ablation
C2985392|T061|argon beam coagulator ablation
C1336817|T191|Transplant-Related Bladder Urothelial Carcinoma
C1336817|T191|Transplant-Related Bladder Transitional Cell Carcinoma
C0855118|T191|Recurrent Follicular Lymphoma
C0855118|T191|Follicle center lymphoma, follicular grade I, II, III recurrent
C0855118|T191|Follicle centre lymphoma, follicular grade I, II, III recurrent
C115384|T191|Recurrent Olfactory Neuroblastoma
C0855020|T191|Recurrent Lentigo Maligna Melanoma
C0855020|T191|Lentigo maligna recurrent
C0855020|T191|Lentigo Maligna Recurrent
C0235813|T191|Neonatal Leukemia
C0235813|T191|LEUKAEMIA NEONATAL
C0235813|T191|Leukaemia neonatal
C0235813|T191|Neonatal leukemia
C0235813|T191|Neonatal leukaemia
C0235813|T191|LEUKEMIA NEONATAL
C0235813|T191|Leukemia neonatal
CL411846|T191|Metastatic Malignant Neoplasm to the Leptomeninges
CL411846|T191|Leptomeningeal Metastasis
CL411846|T191|Leptomeningeal metastases, NOS
CL411846|T191|Leptomeningeal Metastases
CL411846|T191|Metastatic Tumor to the Leptomeninges
CL411846|T191|Metastatic Neoplasm to the Leptomeninges
CL411846|T191|leptomeningeal metastasis
CL411846|T191|Metastasis to the Leptomeninges
CL411846|T191|carcinomatous meningitis
CL411846|T191|meningeal metastasis
CL411846|T191|neoplastic meningitis
CL411846|T191|leptomeningeal carcinoma
C0559185|T191|Adult Spinal Cord Glioblastoma
C0559185|T191|Glioblastoma multiforme of spinal cord (disorder)
C0559185|T191|Glioblastoma multiforme of spinal cord
C0559185|T191|Adult Spinal Cord Glioblastoma Multiforme
C2698751|T191|Pediatric Nodal Marginal Zone Lymphoma
C2698751|T191|Childhood Nodal Marginal Zone Lymphoma
C1300515|T201|Tumor size, invasive component, additional dimension
C1300515|T201|Tumor size, invasive component, additional dimension (observable entity)
C1300515|T201|Tumour size, invasive component, additional dimension
C0008838|T197|Cisplatin
C0008838|T197|DICHLORODIAMMINEPLATINUM CIS 02
C0008838|T197|(SP-4-2)-Diamminedichloroplatinum
C0008838|T197|Cisplatin (substance)
C0008838|T197|cis-platinum
C0008838|T197|cis-Platinum
C0008838|T197|cisplatin
C0008838|T197|Cisplatina
C0008838|T197|(SP-4-2)-diamminedichloroplatinum
C0008838|T197|Cysplatyna
C0008838|T197|119875
C0008838|T197|Diamminodichloride, Platinum
C0008838|T197|PDD
C0008838|T197|Cis-dichloroammine Platinum (II)
C0008838|T197|Platinol-AQ VHA Plus
C0008838|T197|Briplatin
C0008838|T197|cis-Platinum II
C0008838|T197|Metaplatin
C0008838|T197|platinum diamminodichloride
C0008838|T197|Platinum
C0008838|T197|cis-platinum II
C0008838|T197|DDP
C0008838|T197|8041
C0008838|T197|Cis-platinum II Diamine Dichloride
C0008838|T197|Cis-diamminedichloro Platinum (II)
C0008838|T197|Abiplatin
C0008838|T197|Platinum Diamminodichloride
C0008838|T197|Cis-platinum II
C0008838|T197|Cis-diamminedichloridoplatinum
C0008838|T197|platinum, diaminedichloro-, cis- (8CI)
C0008838|T197|cis Platinum
C0008838|T197|cis-diamminedichloro platinum (II)
C0008838|T197|Plastistil
C0008838|T197|Platinol- AQ
C0008838|T197|Platosin
C0008838|T197|Platinum, diamminedichloro-, (SP-4-2)-
C0008838|T197|Citosin
C0008838|T197|Cis-platinum
C0008838|T197|Cis-platinous Diamine Dichloride
C0008838|T197|Cisplatin (product)
C0008838|T197|Platinol-AQ
C0008838|T197|cis-Diamminedichloroplatinum(II)
C0008838|T197|Cis-diammine-dichloroplatinum
C0008838|T197|cis platinum compound
C0008838|T197|DIAMMINEDICHLOROPLATINUM CIS 02
C0008838|T197|Platamine
C0008838|T197|Diaminedichloroplatinum
C0008838|T197|cis-Diaminedichloroplatinum
C0008838|T197|CISplatin
C0008838|T197|Citoplatino
C0008838|T197|CACP
C0008838|T197|Platinoxan
C0008838|T197|CPDD
C0008838|T197|Platistin
C0008838|T197|CDDP
C0008838|T197|Platinex
C0008838|T197|Placis
C0008838|T197|Cismaplat
C0008838|T197|cis dichlorodiammineplatinum
C0008838|T197|cis-platinum II diamine dichloride
C0008838|T197|Platinol
C0008838|T197|cis-Dichlorodiammineplatinum(II)
C0008838|T197|platinol
C0008838|T197|Neoplatin
C0008838|T197|cis-diamminedichloroplatinum
C0008838|T197|Platinum, Diaminedichloro-, cis- (8CI)
C0008838|T197|cis Diamminedichloroplatinum
C0008838|T197|cis-diammine-dichloroplatinum
C0008838|T197|Peyrone's Salt
C0008838|T197|Cisplatyl
C0008838|T197|Peyrone's Chloride
C0008838|T197|cis diamminedichloroplatinum
C0008838|T197|15663-27-1
C0008838|T197|Cisplatin product
C0008838|T197|CDDP - Cisplatin
C0008838|T197|Dichlorodiammineplatinum
C0008838|T197|cis-platinous diamine dichloride
C0008838|T197|Cisplatinum
C0008838|T197|Blastolem
C0008838|T197|Platiblastin
C0008838|T197|cis-Diamminedichloroplatinum
C0008838|T197|Cisplatin [Chemical/Ingredient]
C0008838|T197|Platiblastin-S
C0008838|T197|Lederplatin
C0008838|T197|Platiran
C0008838|T197|cis-Platinum compound
C0008838|T197|cisplatinum
C0008838|T197|cis-DDP
C0008838|T197|Cis-diamminedichloroplatinum
C0008838|T197|CISPLATIN
C0279606|T191|Childhood Hepatocellular Carcinoma
C0279606|T191|Childhood Carcinoma of Liver Cell
C0279606|T191|Childhood Liver Cell Carcinoma
C0279606|T191|Pediatric Carcinoma of the Liver Cell
C0279606|T191|pediatric hepatocellular carcinoma
C0279606|T191|Pediatric Hepatoma
C0279606|T191|hepatoma, childhood
C0279606|T191|Childhood Hepatoma
C0279606|T191|hepatoma, pediatric
C0279606|T191|childhood hepatocellular carcinoma
C0279606|T191|Pediatric Hepatocellular Carcinoma
C0279606|T191|hepatocellular carcinoma, childhood
C0279606|T191|carcinoma, hepatocellular, childhood
C0279606|T191|Pediatric Carcinoma of Liver Cell
C0279606|T191|Pediatric Liver Cell Carcinoma
C0279606|T191|Childhood Carcinoma of the Liver Cell
C0278590|T191|Recurrent Ewing Sarcoma
C0278590|T191|Recurrent Ewing's Sarcoma
C0278590|T191|Ewing's sarcoma recurrent
C0278590|T191|Ewing's tumour recurrent
C0278590|T191|recurrent Ewing's sarcoma
C0278590|T191|Relapsed Ewing's Sarcoma
C0278590|T191|Ewing's sarcoma, recurrent
C0278590|T191|Ewing's Sarcoma, Recurrent
C0278590|T191|Ewing's tumor recurrent
C0280365|T191|Recurrent Oral Cavity Verrucous Carcinoma
C0280365|T191|Relapsed Oral Cavity Verrucous Carcinoma
C0280365|T191|recurrent verrucous carcinoma of the oral cavity
C0280365|T191|verrucous carcinoma of the oral cavity, recurrent
C0280365|T191|Recurrent Verrucous Carcinoma of Mouth
C0280365|T191|Relapsed Verrucous Carcinoma of Oral Cavity
C0280365|T191|Recurrent Verrucous Carcinoma of Oral Cavity
C0280365|T191|Relapsed Verrucous Carcinoma of Mouth
C0280365|T191|Recurrent Verrucous Carcinoma of the Mouth
C0280365|T191|Verrucous carcinoma of the oral cavity recurrent
C0280365|T191|Recurrent Mouth Verrucous Carcinoma
C0280365|T191|oral cavity verrucous carcinoma, recurrent
C0280365|T191|Relapsed Verrucous Carcinoma of the Mouth
C0280365|T191|Relapsed Mouth Verrucous Carcinoma
C0280365|T191|Relapsed Verrucous Carcinoma of the Oral Cavity
C0280365|T191|Recurrent Verrucous Carcinoma of the Oral Cavity
C1332241|T191|Ameloblastic Carcinoma-Secondary Type (Dedifferentiated)
C1332241|T191|Ameloblastic Carcinoma Ex Ameloblastoma
CL448320|T191|Childhood Brain Germ Cell Tumor
CL448320|T191|brain tumor, intracranial germ cell, childhood
CL448320|T191|brain tumor, germ cell, childhood
CL448320|T191|Germ Cell Tumor of Childhood Brain
CL448320|T191|childhood brain tumor, germ cell
CL448320|T191|Germ Cell Neoplasm of the Pediatric Brain
CL448320|T191|childhood brain tumor, intracranial germ cell
CL448320|T191|brain tumor, pediatric, germ cell
CL448320|T191|brain tumor, childhood, germ cell
CL448320|T191|Childhood Brain Germ Cell Neoplasm
CL448320|T191|Germ Cell Neoplasm of Childhood Brain
CL448320|T191|Pediatric Brain Germ Cell Tumor
CL448320|T191|Germ Cell Neoplasm of Pediatric Brain
CL448320|T191|Childhood Germ Cell Brain Tumor
CL448320|T191|Germ Cell Tumor of the Pediatric Brain
CL448320|T191|germ cell brain tumor, childhood
CL448320|T191|childhood germ cell brain tumor
CL448320|T191|intracranial germ cell brain tumor, childhood
CL448320|T191|brain tumor, pediatric, intracranial germ cell
CL448320|T191|Germ Cell Tumor of Pediatric Brain
CL448320|T191|Childhood Germ Cell Brain Neoplasm
CL448320|T191|brain tumor, childhood, intracranial germ cell
CL448320|T191|Pediatric Brain Germ Cell Neoplasm
CL448320|T191|Germ Cell Neoplasm of the Childhood Brain
CL448320|T191|Germ Cell Tumor of the Childhood Brain
C0854797|T191|Resectable Hepatoblastoma
C0854797|T191|Hepatoblastoma, Resectable
C0854797|T191|Hepatoblastoma resectable
C0935681|T191|Non-Hematologic Malignancy
C0935681|T191|nonhematologic cancer
C0935681|T191|Non-Hematologic Cancer
C0853879|T191|Invasive Breast Carcinoma
C0853879|T191|Invasive Carcinoma of Breast
C0853879|T191|Invasive breast carcinoma
C0853879|T191|infiltrating breast cancer
C0853879|T191|Breast Cancer - Invasive
C0853879|T191|Infiltrating Breast Carcinoma
C0853879|T191|Invasive Carcinoma of the Breast
C0853879|T191|invasive breast cancer
C0853879|T191|Breast cancer invasive NOS
C0853879|T191|Infiltrating Carcinoma of the Breast
C0853879|T191|Infiltrating Carcinoma of Breast
C0853879|T191|Invasive Breast Cancer
C2985438|T049|Novel Mutation
C2985438|T049|novel mutation
C1710042|T191|Secondary Osteosarcoma
C1710042|T191|Secondary Bone Osteosarcoma
C0065879|T110|Megestrol Acetate
C0065879|T110|BDH 1298
C0065879|T110|6-Dehydro-6-methyl-17.alpha.-acetoxyprogesterone
C0065879|T110|6-Dehydro-6-methyl-17 alpha-acetoxyprogesterone
C0065879|T110|6-Methyl-6-dehydro-17.alpha.-acetoxyprogesterone
C0065879|T110|(9beta,10alpha)-17-(Acetyloxy)-6-methylpregna-4,6-diene-3,20-dione
C0065879|T110|Maygace
C0065879|T110|Pallace
C0065879|T110|Ovaban
C0065879|T110|17-Hydroxy-6-methylpregna-4,6-diene-3,20-dione acetate
C0065879|T110|Niagestin
C0065879|T110|MEGESTROL ACETATE
C0065879|T110|Megace
C0065879|T110|17 Alpha-acetoxy-6-methylpregna-4,6-diene-3,20-dione
C0065879|T110|BDH-1298
C0065879|T110|Megestil
C0065879|T110|17.alpha.-Acetoxy-6-methylpregna-4,6-diene-3,20-dione
C0065879|T110|Megestat
C0065879|T110|6-Methyl-delta-4,6-pregnadien-17 alpha-ol-3,20-dione Acetate
C0065879|T110|17-Hydroxy-6-methylpregna-4,6-diene-3,20-dione Acetate
C0065879|T110|SC-10363
C1334606|T191|Malignant Neoplasm by Grade
C2698203|T191|Metastatic Ductal Breast Carcinoma
C1377914|T191|Adult Brain Stem Gliosarcoma
C1377914|T191|gliosarcoma, adult brain stem
C1377914|T191|adult brainstem gliosarcoma
C1377914|T191|Adult Brainstem Gliosarcoma
C1377914|T191|gliosarcoma, adult brainstem
C1377914|T191|adult brain stem gliosarcoma
C0278811|T191|Unresectable Extrahepatic Bile Duct Carcinoma
C0278811|T191|Unresectable Cancer of the Extrahepatic Bile Duct
C0278811|T191|Unresectable Extrahepatic Bile Duct Cancer
C0278811|T191|unresectable extrahepatic bile duct cancer
C0278811|T191|Non-Resectable Extrahepatic Bile Duct Carcinoma
C0278811|T191|Unresectable Cancer of Extrahepatic Bile Duct
C0278811|T191|bile duct cancer, unresectable extrahepatic
C0278811|T191|extrahepatic bile duct cancer, unresectable
C0541315|T121|Everolimus
C0541315|T121|42-O-(2-hydroxy)ethyl rapamycin
C0541315|T121|42-O-(2-Hydroxy)ethyl Rapamycin
C0541315|T121|SDZ-RAD
C0541315|T121|(1R,9S,12S,15R,16E,18R,19R,21R,23S,24E,26E,28E,30S,32S,35R)-1,18-Dihydroxy-12-((1R)-2-((1S,3R,4R)-4-(2-hydroxyethoxy)-3-methoxycyclohexyl)-1-methylethyl)-19,30-dimethoxy-15,17,21,23,29,35-hexamethyl-11,36-dioxa-4-azatricyclo(30.3.1.04,9)hexatriaconta-16,24,26,28-tetraene-2,3,10,14,20-pentaone
C0541315|T121|EVEROLIMUS
C0541315|T121|40-O-(2-hydroxyethyl)-rapamycin
C0541315|T121|Afinitor
C0541315|T121|Everolimus (product)
C0541315|T121|RAD 001
C0541315|T121|RAD001
C0541315|T121|Certican
C0541315|T121|SDZ RAD
C0541315|T121|Everolimus (substance)
C0541315|T121|everolimus
C0279556|T191|Invasive Ductal Breast Carcinoma with Predominant Intraductal Component
C0279556|T191|Infiltrating Ductal Breast Carcinoma with Predominant Intraductal Component
C1709352|T033|Ossified Mass
C0445036|T033|M1a Stage Finding
C0445036|T033|M1a Stage
C0445036|T033|M1a TNM Finding
C0445036|T033|Metastasis stage M1a (finding)
C0445036|T033|M1a Metastasis Finding
C0445036|T033|Metastasis stage M1a
C0445036|T033|M1a Distant Metastasis Stage Finding
C0445036|T033|M1a Cancer Stage Finding
C0445036|T033|M1a Distant Metastasis Finding
C0445036|T033|Metastasis Stage M1a
C0445036|T033|M1a Metastasis Stage
C0445036|T033|M1a
C0153677|T191|Metastatic Malignant Neoplasm to the Mediastinum
C0153677|T191|Metastatic Neoplasm to the Mediastinum
C0153677|T191|Metastases to Mediastinum
C0153677|T191|Metastasis to the Mediastinum
C0153677|T191|Metastatic Tumor to the Mediastinum
C0153677|T191|Metastases to the Mediastinum
C3273727|T191|Breast Solid Neuroendocrine Carcinoma
C0854779|T191|Recurrent Rectosigmoid Carcinoma
C0854779|T191|Rectosigmoid Cancer, Recurrent
C0854779|T191|Relapsed Rectosigmoid Cancer
C0854779|T191|Recurrent Rectosigmoid Cancer
C0854779|T191|Rectosigmoid cancer recurrent
C0278736|T191|Stage II Childhood Lymphoblastic Lymphoma
C0278736|T191|Pediatric Lymphoblastic Lymphoma Stage II
C0278736|T191|Childhood Lymphoblastic Lymphoma Stage II
C0278736|T191|Stage II Pediatric Lymphoblastic Lymphoma
C0278736|T191|Stage II Childhood Precursor Lymphoblastic Lymphoma
C0279603|T191|Chondroblastic Osteosarcoma
C0279603|T191|Chondroblastic osteosarcoma (morphologic abnormality)
C0279603|T191|osteosarcoma, chondroblastic
C0279603|T191|chondroblastic osteosarcoma
C0279603|T191|chondrosarcomatous osteogenic sarcoma
C0279603|T191|Chondroblastic Osteogenic Sarcoma
C0279603|T191|osteogenic sarcoma, chondrosarcomatous
C0279603|T191|chondroblastic osteogenic sarcoma
C0279603|T191|osteogenic sarcoma, chondroblastic
C0279603|T191|chondrosarcomatous osteosarcoma
C0279603|T191|Chondroblastic osteosarcoma
C0279603|T191|Osteochondrosarcoma
C0279603|T191|Chondrosarcomatous osteosarcoma
C0279603|T191|osteosarcoma, chondrosarcomatous
C0279603|T191|sarcoma, osteogenic, chondrosarcomatous
C0334579|T191|Anaplastic Astrocytoma
C0334579|T191|anaplastic astrocytoma
C0334579|T191|Astrocytoma, anaplastic
C0334579|T191|Grade III Astrocytoma
C0334579|T191|GRADE III ASTROCYTOMA
C0334579|T191|astrocytoma WHO grade III
C0334579|T191|ASTROCYTOMA, ANAPLASTIC, MALIGNANT
C0334579|T191|Malignant astrocytoma
C0334579|T191|GRADE III ASTROCYTIC TUMOR
C0334579|T191|Grade III Astrocytic Tumor
C0334579|T191|Grade III Astrocytomas
C0334579|T191|MALIGNANT ASTROCYTOMA
C0334579|T191|Astrocytoma, Grade III
C0334579|T191|Anaplastic Astrocytomas
C0334579|T191|Astrocytomas, Anaplastic
C0334579|T191|Astrocytoma, Anaplastic
C0334579|T191|Astrocytoma malignant
C0334579|T191|Anaplastic astrocytoma
C0334579|T191|Astrocytomas, Grade III
C0334579|T191|Malignant Astrocytoma
C0334579|T191|Grade III Astrocytic Neoplasm
C0334579|T191|Astrocytoma malignant NOS
C0334579|T191|Astrocytoma, anaplastic (morphologic abnormality)
C0334579|T191|GRADE III ASTROCYTIC NEOPLASM
C1334273|T191|Invasive Breast Carcinoma by Histologic Grade
C1334273|T191|Infiltrating Breast Carcinoma by Histologic Grade
C1334273|T191|Infiltrating Breast Carcinoma by Nottingham Combined Histologic Grade
C1334273|T191|Invasive Breast Carcinoma by Nottingham Combined Histologic Grade
C0700476|T116|Goserelin Acetate
C0700476|T116|ZDX
C0700476|T116|Acetate, Goserelin
C0700476|T116|goserelin acetate
C0700476|T116|Goserelin acetate preparation
C0700476|T116|Goserelin Acetate [Chemical/Ingredient]
C0700476|T116|Goserelin acetate preparation (product)
C0700476|T116|D-Ser(bu(t))(6)azgly(10)-LHRH Acetate
C0700476|T116|Goserelin acetate (substance)
C0700476|T116|GOSERELIN ACETATE
C0700476|T116|Goserelin acetate
C0700476|T116|Zoladex
C0280096|T191|Adenocarcinoma of Unknown Primary
C0854750|T191|Recurrent Colorectal Carcinoma
C0854750|T191|Colorectal Cancer, Recurrent
C0854750|T191|Colorectal cancer recurrent
C0854750|T191|Colorectal Carcinoma Recurrent
C0854750|T191|Recurrent Colorectal Cancer
CL448706|T045|Targeted Mutation
CL448706|T045|Targeted Modification
CL448706|T045|Targeted DNA Alteration
CL448706|T045|Targeted Sequence Alteration
CL448706|T045|Targeted DNA Modification
C1709664|T191|Primary Intraosseous Squamous Cell Carcinoma Derived From Keratocystic Odontogenic Tumor
C1709664|T191|Primary Intraosseous Carcinoma Ex Keratocystic Odontogenic Tumor
C1273120|T033|Polyp size, additional dimension
C1273120|T033|Polyp size, additional dimension (observable entity)
C1273120|T033|Polyp size additional dimensions
C1334723|T191|Metastatic Malignant Neoplasm to the Adult Brain
C1334723|T191|Metastasis to the Adult Brain
C1334723|T191|Metastatic Tumor to the Adult Brain
C1334723|T191|Brain Metastases, Adult
C1334723|T191|Metastatic Neoplasm to the Adult Brain
C1334723|T191|Secondary Malignant Neoplasm to the Adult Brain
C1334723|T191|Secondary Malignant Tumor to the Adult Brain
C1335760|T033|Resectable Mass
C1335760|T033|Resected Mass
C0854769|T191|Recurrent Esophageal Squamous Cell Carcinoma
C0854769|T191|Oesophageal squamous cell carcinoma recurrent
C0854769|T191|Recurrent Squamous Cell Carcinoma of Esophagus
C0854769|T191|Oesophageal squamous cell carcinoma site unspecified recurrent
C0854769|T191|Recurrent Squamous Cell Carcinoma of the Esophagus
C0854769|T191|Esophageal squamous cell carcinoma site unspecified recurrent
C0854769|T191|Esophageal squamous cell carcinoma recurrent
C0281700|T191|Stage I Childhood Burkitt Lymphoma
C0281700|T191|Stage I Pediatric Small Non-Cleaved Cell Lymphoma
C0281700|T191|Childhood Small Non-Cleaved Cell Lymphoma Stage I
C0281700|T191|Stage I Childhood Small Non-Cleaved Cell Lymphoma
C0281700|T191|Pediatric Small Non-Cleaved Cell Lymphoma Stage I
C0281700|T191|Stage I Childhood Burkitt's Lymphoma
C1708397|T191|Hydroa Vacciniforme-Like Lymphoma
C1708397|T191|Hydroa Vacciniforme-Like Cutaneous T-Cell Lymphoma
C0854909|T191|Anaplastic (Malignant) Intracranial Meningioma
C535837|T191|Hereditary Pancreatic Carcinoma
C535837|T191|Familial Pancreatic carcinoma
C535837|T191|Familial Pancreatic Cancer
C535837|T191|pancreatic cancer, familial
C535837|T191|Familial Pancreatic Carcinoma
C535837|T191|Hereditary Pancreatic Cancer
C535837|T191|Pancreatic carcinoma, familial
C535837|T191|familial pancreatic cancer
C535837|T191|hereditary pancreatic cancer
C535837|T191|pancreatic cancer, hereditary
C1335460|T191|Postsurgical Stage IV Hepatoblastoma
C1512224|T191|Glycogen-Rich, Clear Cell Breast Carcinoma
C1513365|T191|Mixed Epithelial/Mesenchymal Metaplastic Breast Carcinoma
C1513365|T191|Breast Carcinosarcoma
C1334798|T191|Monomorphic Post-Transplant Lymphoproliferative Disorder
C1334798|T191|Post-transplant lymphoproliferative disorder (Monoclonal), NOS
C1334798|T191|PTLD (Monoclonal)
C1334798|T191|Monomorphic PTLD
C1300514|T201|Tumor size, invasive component, greatest dimension
C1300514|T201|Tumour size, invasive component, greatest dimension
C1300514|T201|Tumor size, invasive component, greatest dimension (observable entity)
C1709093|T049|Multiple Transition Abnormalities
C1709093|T049|Multiple Transition Mutations
C1709093|T049|Transition Mutations
C1333991|T191|Lynch 2 Syndrome
C1333991|T191|Colorectal Cancer, Hereditary Nonpolyposis, Type 2
C1333991|T191|COLON CANCER, FAMILIAL NONPOLYPOSIS, TYPE 2
C1333991|T191|COLORECTAL CANCER, HEREDITARY NONPOLYPOSIS, TYPE 2
C1333991|T191|Lynch Syndrome II [Disease/Finding]
C1333991|T191|Lynch Cancer Family Syndrome II
C1333991|T191|LYNCH SYNDROME II
C1333991|T191|COCA2
C1333991|T191|Lynch Syndrome II
C1333991|T191|FCC2
C1333991|T191|Colon Cancer, Familial Nonpolyposis, Type 2
C1333991|T191|HNPCC2
C1333991|T191|Familial Non-Polyposis Colon Cancer Type 2
C1333991|T191|Hereditary Non-Polyposis Colon Cancer Type 2
C1332964|T191|Childhood Clear Cell Sarcoma of Soft Parts
C1332964|T191|Pediatric Clear Cell Sarcoma of Soft Parts
C0280427|T191|Recurrent Adult T-Cell Leukemia/Lymphoma
C0280427|T191|Recurrent HTLV-1 Associated Adult T-Cell Lymphoma/Leukemia
C0280427|T191|Adult T-Cell Lymphoma/Leukemia Recurrent
C0280427|T191|Recurrent Adult T-Cell Lymphoma/Leukemia
C0280427|T191|HTLV-1 Associated Adult T-Cell Lymphoma/Leukemia Relapsed
C0280427|T191|Relapsed HTLV-1 Associated Adult T-Cell Lymphoma/Leukemia
C0280427|T191|HTLV-1 Associated Adult T-Cell Lymphoma/Leukemia Recurrent
C1512746|T191|Infiltrating Bladder Urothelial Carcinoma with Giant Cells
C1265601|T190|Solitary Mass
C1265601|T190|Solitary mass
C1265601|T190|Single mass
C1265601|T190|Solitary mass (morphologic abnormality)
C1541317|T191|Adult Gliosarcoma
C1541317|T191|adult gliosarcoma
C1541317|T191|gliosarcoma, adult
CL448337|T191|Stage I Bladder Urothelial Carcinoma
CL448337|T191|Stage I Transitional Cell Carcinoma of Urinary Bladder
CL448337|T191|Stage I Urinary Bladder Transitional Cell Carcinoma
CL448337|T191|Stage I Transitional Cell Carcinoma of the Urinary Bladder
CL448337|T191|Stage I Bladder Urothelial Carcinoma AJCC v6
CL448337|T191|Stage I Bladder Urothelial Carcinoma AJCC v7
CL448337|T191|Stage I Transitional Cell Carcinoma of the Bladder
CL448337|T191|Stage I Transitional Cell Carcinoma of Bladder
C1518362|T061|Radiation, Non-Ionizing DX or RX
C0162735|T045|Point Mutation
C0162735|T045|Mutation, Point
C0162735|T045|Mutations, Point
C0162735|T045|point mutation
C0162735|T045|Point Mutations
C0162735|T045|Point mutation (finding)
C0162735|T045|Point mutation
C0347021|T191|Metastatic Malignant Neoplasm to the Choroid
C0347021|T191|Metastatic Tumor to the Choroid
C0347021|T191|Metastatic Neoplasm to the Choroid
C0153685|T191|Metastatic Malignant Neoplasm to the Kidney
C0153685|T191|Metastasis to Kidney
C0153685|T191|Metastases to the Kidney
C0153685|T191|Metastatic Neoplasm to the Kidney
C0153685|T191|Renal Metastasis
C0153685|T191|Metastasis to the Kidney
C0153685|T191|Renal Metastases
C0153685|T191|Metastatic Tumor to the Kidney
C0153685|T191|Metastases to Kidney
C0877294|T191|Metastatic Malignant Neoplasm to the Placenta
C0877294|T191|Metastasis to the Placenta
C0877294|T191|Metastasis to Placenta
C0877294|T191|Metastatic Tumor to the Placenta
C0877294|T191|Metastatic Neoplasm to the Placenta
C0854822|T191|Stage I Anaplastic Large Cell Lymphoma
C0854822|T191|Anaplastic Large Cell Lymphoma T- and Null-Cell Types Stage I
C0854822|T191|Anaplastic Large Cell Lymphoma Stage I
C0279942|T191|Metastatic Childhood Soft Tissue Sarcoma
C0279942|T191|Metastatic Childhood Sarcoma of Soft Tissue
C0279942|T191|Metastatic Pediatric Sarcoma of the Soft Tissue
C0279942|T191|pediatric metastatic STS
C0279942|T191|soft tissue sarcoma, childhood, metastatic
C0279942|T191|Metastatic Childhood Sarcoma of the Soft Tissue
C0279942|T191|STS, metastatic, childhood
C0279942|T191|childhood STS, metastatic
C0279942|T191|pediatric STS, metastatic
C0279942|T191|metastatic childhood soft tissue sarcoma
C0279942|T191|childhood soft tissue sarcoma, metastatic
C0279942|T191|childhood metastatic STS
C0279942|T191|Metastatic Pediatric Soft Tissue Sarcoma
C0279942|T191|Metastatic Pediatric Sarcoma of Soft Tissue
C0686068|T191|Metastatic Malignant Neoplasm to the Stomach
C1332997|T191|Childhood T Lymphoblastic Leukemia/Lymphoma
C1332997|T191|Childhood Precursor T-Lymphoblastic Lymphoma/Leukemia
C0278530|T191|Recurrent Adult Hodgkin Lymphoma
C0278530|T191|HD, adult, relapsed
C0278530|T191|relapsed adult HD
C0278530|T191|HD, recurrent, adult
C0278530|T191|Hodgkin's lymphoma, relapsed, adult
C0278530|T191|recurrent adult Hodgkin's disease
C0278530|T191|Recurrent Adult Hodgkin's Lymphoma
C0278530|T191|adult Hodgkin's disease, recurrent
C0278530|T191|adult HD, relapsed
C0278530|T191|relapsed adult Hodgkin's disease
C0278530|T191|relapsed Hodgkin's disease, adult
C0278530|T191|adult Hodgkin's disease, relapsed
C0278530|T191|adult HD, recurrent
C0278530|T191|recurrent HD, adult
C0278530|T191|recurrent adult HD
C0278530|T191|HD, adult, recurrent
C0278530|T191|recurrent adult Hodgkin lymphoma
C0278530|T191|Hodgkin's disease, relapsed, adult
C0278530|T191|Relapsed Adult Hodgkin's Lymphoma
C0278530|T191|lymphoma, relapsed adult Hodgkin's
C0278530|T191|Recurrent Adult Hodgkin's Disease
C0278530|T191|Relapsed Adult Hodgkin's Disease
C0278530|T191|recurrent Hodgkin's disease, adult
C0278530|T191|HD, relapsed, adult
C1332055|T191|AIDS-Related Plasmablastic Lymphoma
C0854983|T191|Recurrent Lung Adenocarcinoma
C0854983|T191|Recurrent Adenocarcinoma of Lung
C0854983|T191|Lung adenocarcinoma recurrent
C0854983|T191|Adenocarcinoma of lung recurrent
C0854983|T191|Lung Adenocarcinoma, Recurrent
C0854983|T191|Recurrent Adenocarcinoma of the Lung
C2986686|T191|Stage IV AIDS-Related Lymphoma
C2986686|T191|stage IV AIDS-related lymphoma
C0023452|T191|Childhood Acute Lymphoblastic Leukemia
C0023452|T191|childhood ALL
C0023452|T191|pediatric ALL
C0023452|T191|Acute lymphocytic leukemia (ALL), child
C0023452|T191|Childhood Precursor Lymphoblastic Leukemia
C0023452|T191|Childhood Acute Lymphoid Leukemia
C0023452|T191|L1 Lymphocytic Leukemia
C0023452|T191|Leukemia, Lymphocytic, Acute, L1
C0023452|T191|Leukemia, Lymphoblastic, Acute, L1
C0023452|T191|Leukemia, L1 Lymphocytic
C0023452|T191|pediatric acute lymphoblastic leukemia
C0023452|T191|leukemia, acute lymphoblastic, pediatric
C0023452|T191|pediatric acute lymphogenous leukemia
C0023452|T191|childhood precursor lymphoblastic leukemia
C0023452|T191|Pediatric Acute Lymphoid Leukemia
C0023452|T191|lymphoblastic leukemia, acute, childhood
C0023452|T191|pediatric acute lymphoid leukemia
C0023452|T191|childhood acute lymphoblastic leukemia
C0023452|T191|leukemia, acute lymphoblastic, childhood
C0023452|T191|ALL, Childhood
C0023452|T191|Childhood Acute Lymphocytic Leukemia
C0023452|T191|ALL, pediatric
C0023452|T191|ALL, childhood
C0023452|T191|lymphoblastic leukemia, acute, pediatric
C0023452|T191|Pediatric ALL
C0023452|T191|Lymphocytic Leukemia, L1
C0023452|T191|childhood acute lymphoid leukemia
C0023452|T191|Pediatric Acute Lymphocytic Leukemia
C0023452|T191|childhood leukemia, acute lymphoblastic
C0023452|T191|Childhood ALL
C0023452|T191|acute lymphoblastic leukemia, pediatric
C0023452|T191|childhood acute lymphocytic leukemia
C0023452|T191|Lymphoblastic Leukemia, Acute, L1
C0023452|T191|childhood acute lymphogenous leukemia
C0023452|T191|Childhood Acute Lymphogenous Leukemia
C0023452|T191|Leukemia, acute lymphocytic (ALL), child
C0023452|T191|Lymphoblastic Leukemia, Acute, Childhood
C0023452|T191|Pediatric Acute Lymphoblastic Leukemia
C0023452|T191|Pediatric Acute Lymphogenous Leukemia
C0023452|T191|acute lymphoblastic leukemia, childhood
C0023452|T191|Pediatric Acute Lymphocytic Leukemia (ALL)
C0023452|T191|pediatric acute lymphocytic leukemia
C1335964|T191|Signet Ring Cell Breast Carcinoma
C1335964|T191|Primary Signet Ring Cell Carcinoma of the Breast
C1335964|T191|SRC Carcinoma of Breast
C1335964|T191|SRC Carcinoma of the Breast
C1335964|T191|Signet Ring Cell Carcinoma of the Breast
C1335964|T191|Primary SRC Breast Carcinoma
C1335964|T191|Primary Signet Ring Cell Carcinoma of Breast
C1335964|T191|Signet Ring Cell Carcinoma of Breast
C1335964|T191|Mammary Signet Ring Cell Carcinoma
C1335964|T191|Primary Signet Ring Cell Breast Carcinoma
C1335964|T191|Primary SRC Carcinoma of the Breast
C1335964|T191|Primary SRC Carcinoma of Breast
C1335964|T191|Primary Mammary Signet Ring Cell Carcinoma
C1335964|T191|SRC Breast Carcinoma
C0677922|T061|Ovarian Ablation
C0677922|T061|ovarian suppression
C0677922|T061|ovarian ablation
C0677922|T061|Ovarian ablation
C0677922|T061|Ovarian ablation (procedure)
C1709018|T033|Microcalcification Present in Neoplastic and Non-Neoplastic Tissue
C0241353|T033|Testicular Mass
C0241353|T033|Testicular lump
C0241353|T033|Mass of testis
C0241353|T033|TESTICULAR MASS
C0241353|T033|TESTES MASS
C0241353|T033|Mass of testicle
C0241353|T033|TESTIS MASS
C0241353|T033|Mass of testicle (finding)
C0241353|T033|Lump in testis
C0241353|T033|Testicular mass
C1883538|T061|Vinorelbine-Epirubicin Regimen
C1517527|T033|Geographic Necrosis
C1512741|T191|Infiltrating Bladder Urothelial Carcinoma, Nested Variant
C0454270|T081|High-Dose Rate Brachytherapy
C1333420|T191|Epithelial Predominant Pulmonary Blastoma
C0599155|T045|Missense Mutation
C0599155|T045|Non-Synonymous Mutation
C0599155|T045|Substitution Mutation
C0599155|T045|missense mutation
C0599155|T045|Exonic Non-Synonymous Mutation
C0599155|T045|Missense Mutations
C0599155|T045|Exon Non-Synonymous Mutation
C0599155|T045|Mutation, Missense
C0599155|T045|Missense Mutation Abnormality
C0599155|T045|Mutations, Missense
CL449192|T033|N4 Stage Finding
CL472690|T191|Childhood Cerebellar Anaplastic Astrocytoma
CL448305|T191|Recurrent Pharyngeal Carcinoma
CL448305|T191|Recurrent Pharynx Carcinoma
CL448305|T191|Recurrent Pharyngeal Cancer
CL448305|T191|Recurrent Carcinoma of Pharynx
CL448305|T191|Recurrent Cancer of Pharynx
CL448305|T191|Relapsed Pharyngeal Carcinoma
CL448305|T191|Relapsed Carcinoma of Pharynx
CL448305|T191|Recurrent Pharynx Cancer
CL448305|T191|Relapsed Pharyngeal Cancer
CL448305|T191|Pharyngeal Cancer, Recurrent
CL448305|T191|Relapsed Cancer of the Pharynx
CL448305|T191|Relapsed Pharynx Carcinoma
CL448305|T191|Relapsed Pharynx Cancer
CL448305|T191|Relapsed Carcinoma of the Pharynx
CL448305|T191|Relapsed Cancer of Pharynx
CL448305|T191|Recurrent Cancer of the Pharynx
CL448305|T191|Recurrent Carcinoma of the Pharynx
C0278584|T191|Metastatic Carcinoma to the Uterine Cervix
C0278584|T191|Secondary Carcinoma to the Uterine Cervix
C0278584|T191|Metastatic Carcinoma to the Cervix Uteri
C0278584|T191|Metastatic Carcinoma to the Cervix
C0278584|T191|Secondary Carcinoma to the Cervix
C0278584|T191|Secondary Carcinoma to the Cervix Uteri
C1519207|T191|Sebaceous Breast Carcinoma
C1336808|T191|Transplant-Related Carcinoma
C1708566|T191|Invasive Prostate Carcinoma
C1708566|T191|Infiltrating Prostate Carcinoma
C0856022|T191|Recurrent Splenic Marginal Zone Lymphoma
C0856022|T191|Relapsed Splenic Marginal Zone Lymphoma
C0856022|T191|Splenic marginal zone lymphoma recurrent
C0856022|T191|Recurrent Splenic Marginal Zone B-Cell Lymphoma
C1709107|T033|N1c Stage Finding
C1709107|T033|N1c
C1709107|T033|Node Stage N1c
C1709107|T033|N1c Lymph Node Stage
C1709107|T033|N1c TNM Finding
C1709107|T033|N1c Cancer Stage Finding
C1709107|T033|N1c Regional Lymph Node Stage Finding
C1709107|T033|N1c Regional Lymph Nodes Finding
C1709107|T033|N1c Node Stage
C1709107|T033|N1c Lymph Node Finding
C1709107|T033|N1c Stage
C1709107|T033|Lymph Node Stage N1c
C1709107|T033|N1c Node Finding
C0229985|T023|Surgical Margin
C0229985|T023|Surgical margins (body structure)
C0229985|T023|Surgical margins
C0229985|T023|Surgical Margins
C0229985|T023|margin
C0229985|T023|Margins of excision
C3273218|T191|Invasive Lobular Breast Carcinoma, Tubulolobular Variant
CL322961|T169|Apoptosis
CL322961|T169|Gene-directed cell death
CL322961|T169|Programmed Cell Death, Type I
CL322961|T169|programmed cell death by apoptosis
CL322961|T169|type I programmed cell death
CL322961|T169|apoptosis
CL322961|T169|Apoptosis Pathway
CL322961|T169|apoptotic programmed cell death
CL322961|T169|Programmed Cell Death
CL322961|T169|apoptotic process
CL322961|T169|apoptotic cell death
CL322961|T169|Apoptosis (morphologic abnormality)
CL322961|T169|Apoptotic Process
CL322961|T169|programmed cell death
CL322961|T169|PCD
C1848888|T033|Painless Testicular Mass
C1848888|T033|Painless testicular mass
C1333832|T191|Grade 1 Invasive Breast Carcinoma
C1333832|T191|Well Differentiated Invasive Breast Carcinoma
C1333832|T191|Low Combined Histologic Grade Infiltrating Breast Carcinoma
C1333832|T191|Grade 1 Infiltrating Breast Carcinoma
C1333832|T191|Favorable Infiltrating Breast Carcinoma
C1333832|T191|Well Differentiated Infiltrating Breast Carcinoma
C0854917|T191|Rhabdoid Tumor of the Kidney
C0854917|T191|Rhabdoid Neoplasm of the Kidney
C0854917|T191|Rhabdoid tumor of the kidney
C0854917|T191|Malignant Rhabdoid Tumor of Kidney
C0854917|T191|MRTK
C0854917|T191|Rhabdoid Tumor of the Kidney (RTK)
C0854917|T191|Rhabdoid Neoplasm of Kidney
C0854917|T191|Kidney Rhabdoid Tumor
C0854917|T191|Malignant Rhabdoid Tumor of the Kidney
C0854917|T191|Renal Rhabdoid Tumor
C0854917|T191|Renal Rhabdoid Neoplasm
C0854917|T191|Rhabdoid Tumour of Kidney
C0854917|T191|Rhabdoid Tumour of the Kidney
C1882250|T061|PCH Regimen
C1882250|T061|Paclitaxel-Carboplatin-Herceptin Regimen
C1335939|T191|Metastatic Lymphoma to the Heart
C1335939|T191|Secondary Cardiac Lymphoma
C1335939|T191|Secondary Heart Lymphoma
C1708109|T033|Fungating Mass
C1708109|T033|fungating lesion
C1332544|T191|Benzene-Related Acute Myeloid Leukemia
C1332980|T191|Childhood Mature T- and NK-Cell Lymphoma
C1332980|T191|Pediatric Peripheral T Cell Lymphoma
C1332980|T191|Childhood Peripheral T Cell Lymphoma
C0684964|T191|Metastatic Malignant Neoplasm to the Hypopharynx
C0684964|T191|Metastatic Tumor to the Hypopharynx
C0684964|T191|Metastatic Neoplasm to the Hypopharynx
C1708350|T191|Hereditary Leiomyomatosis and Renal Cell Cancer
C1708350|T191|HLRCC
C1708350|T191|Hereditary Leiomyomatosis and Renal Cell Carcinoma
C1708350|T191|hereditary leiomyomatosis and renal cell cancer syndrome
C0278579|T191|Recurrent Cervical Carcinoma
C0278579|T191|recurrent cervix cancer
C0278579|T191|Relapsed Cervix Carcinoma
C0278579|T191|carcinoma of the cervix, recurrent
C0278579|T191|Cervical Carcinoma Recurrent
C0278579|T191|Recurrent Carcinoma of Cervix
C0278579|T191|Recurrent Carcinoma of Uterine Cervix
C0278579|T191|Relapsed Carcinoma of the Cervix Uteri
C0278579|T191|Relapsed Cervical Carcinoma
C0278579|T191|Carcinoma cervix recurrent
C0278579|T191|uterine cervical cancer, recurrent
C0278579|T191|recurrent cervical cancer
C0278579|T191|Relapsed Carcinoma of the Uterine Cervix
C0278579|T191|Relapsed Carcinoma of Cervix
C0278579|T191|Relapsed Cervix Uteri Carcinoma
C0278579|T191|Recurrent Carcinoma of the Cervix
C0278579|T191|cervix cancer recurrent
C0278579|T191|Relapsed Uterine Cervix Carcinoma
C0278579|T191|Relapsed Carcinoma of the Cervix
C0278579|T191|Recurrent Carcinoma of Cervix Uteri
C0278579|T191|Relapsed Carcinoma of Cervix Uteri
C0278579|T191|recurrent carcinoma of the cervix
C0278579|T191|Recurrent Uterine Cervix Carcinoma
C0278579|T191|recurrent cancer of the cervix
C0278579|T191|Relapsed Carcinoma of Uterine Cervix
C0278579|T191|Carcinoma uterine cervix recurrent
C0278579|T191|uterine cervix cancer, recurrent
C0278579|T191|Recurrent Cervix Uteri Carcinoma
C0278579|T191|Cervix carcinoma recurrent
C0278579|T191|Recurrent Carcinoma of the Uterine Cervix
C0278579|T191|cancer of the cervix, recurrent
C0278579|T191|Recurrent Carcinoma of the Cervix Uteri
C0278579|T191|recurrent uterine cervix cancer
C0278579|T191|cervical cancer, recurrent
C0278579|T191|Cervical carcinoma recurrent
C0278579|T191|Recurrent Cervical Cancer
C0278579|T191|Cervical cancer recurrent
C0278579|T191|Cervix uteri cancer recurrent
C1335487|T191|Primary Intraosseous Squamous Cell Carcinoma Derived From Odontogenic Cyst
C1335487|T191|Primary Intraosseous Carcinoma Ex Odontogenic Cyst
C1710670|T061|Whole-Abdominal Irradiation
C0600558|T061|Neoadjuvant Therapy
C0600558|T061|Treatments, Neoadjuvant
C0600558|T061|Neoadjuvant therapy
C0600558|T061|Neoadjuvant Therapies
C0600558|T061|Neoadjuvant Treatments
C0600558|T061|Therapy, Neoadjuvant
C0600558|T061|Preoperative Therapy
C0600558|T061|Induction Therapy
C0600558|T061|Neoadjuvant
C0600558|T061|induction therapy
C0600558|T061|Therapies, Neoadjuvant
C0600558|T061|neoadjuvant therapy
C0600558|T061|Neoadjuvant Treatment
C0600558|T061|Treatment, Neoadjuvant
C0861876|T191|Recurrent Liver Carcinoma
C0861876|T191|Liver, cancer of, recurrent
C0861876|T191|Relapsed Liver Cancer
C0861876|T191|Liver carcinoma recurrent
C0861876|T191|Relapsed Cancer of Liver
C0861876|T191|Carcinoma liver recurrent
C0861876|T191|Relapsed Cancer of the Liver
C0861876|T191|Liver cell carcinoma recurrent
C0861876|T191|Relapsed Hepatic Cancer
C0861876|T191|Recurrent Cancer of Liver
C0861876|T191|Recurrent Cancer of the Liver
C0861876|T191|Recurrent Hepatic Cancer
C0861876|T191|Recurrent Liver Cancer
C0861876|T191|Hepatic cancer recurrent
C1881250|T045|Intronic Mutation
C1881250|T045|Intron Mutation
C1709017|T033|Microcalcification Present in Neoplastic Tissue
C1335937|T191|Metastatic Hodgkin Lymphoma to Cerebral Hemisphere
C1335937|T191|Secondary Cerebral Hodgkin's Lymphoma
C1335937|T191|Secondary Cerebral Hodgkin Lymphoma
C1335937|T191|Secondary Cerebral Hodgkin's Disease
C1335937|T191|Metastatic Hodgkin's Lymphoma to Cerebral Hemisphere
C0686477|T191|Metastatic Malignant Neoplasm to the Retina
C0686477|T191|Metastasis to the Retina
C0686477|T191|Metastatic Neoplasm to the Retina
C0686477|T191|Metastatic Tumor to the Retina
C1333848|T191|Grade 3a Malignant Neoplasm
C0000734|T033|Abdominal Mass
C0000734|T033|Abdominal mass NOS
C0000734|T033|Mass of abdominal cavity structure
C0000734|T033|Abdominal lump
C0000734|T033|Mass in abdomen
C0000734|T033|Abdominal mass
C0000734|T033|Abdominal mass (finding)
C0000734|T033|Intra-abdominal mass
C0000734|T033|Mass of abdominal cavity structure (finding)
C0000734|T033|ABDOMINAL MASS
C1272628|T033|Microcalcification Present in Non-Neoplastic Tissue
C1300693|T201|Lesion size, additional dimension
C1300693|T201|Lesion size, additional dimension (observable entity)
C0854868|T191|Transformed Recurrent Non-Hodgkin Lymphoma
C0854868|T191|NonHodgkin's Lymphoma Transformed Recurrent
C0854868|T191|Non-Hodgkin's Lymphoma Transformed Recurrent
C0854868|T191|Transformed Recurrent Non-Hodgkin's Lymphoma
C1335981|T191|Small Cell Undifferentiated Hepatoblastoma
C0686106|T191|Metastatic Malignant Neoplasm to the Anus
C0686106|T191|Metastatic Malignant Tumor to the Anus
C0079172|T061|Cranial Irradiation
C0079172|T061|Cranial Irradiations
C0079172|T061|Irradiations, Cranial
C0079172|T061|Irradiation, Cranial
C017039|T110|Azastene
C017039|T110|4,4,17-alpha-trimethylandrost-5-eno[2,3,-d]isoxazol-17-ol
C017039|T110|(17 beta)-4,4,17-trimethylandrosta-2,5-diene(3,2-d)isoxazol-17-ol
C017039|T110|isoxazol
C017039|T110|azastene
C017039|T110|AZASTENE
C0346151|T191|Scirrhous Breast Carcinoma
C0346151|T191|Infiltrating Carcinoma of Breast with Fibrotic Stroma
C0346151|T191|Infiltrating Carcinoma of the Breast with Fibrotic Stroma
C0346151|T191|Scirrhous Carcinoma of the Breast
C0346151|T191|Scirrhous Carcinoma of Breast
C0346151|T191|Scirrhous carcinoma of breast
C0346151|T191|Scirrhous carcinoma of breast (disorder)
C0022790|T191|Krukenberg Tumor
C0022790|T191|Krukenberg Tumor [Disease/Finding]
C0022790|T191|Second malig neo ovary
C0022790|T191|Carcinoma, Krukenberg
C0022790|T191|Krukenberg's Tumor
C0022790|T191|Krukenberg Carcinoma
C0022790|T191|Krukenberg Neoplasm
C0022790|T191|Tumor, Krukenberg
C0022790|T191|Krukenburg tumor
C0022790|T191|Secondary malignant neoplasm of ovary
C0022790|T191|Krukenberg tumor
C0022790|T191|Krukenburg tumour
C0022790|T191|Krukenberg tumour
C0022790|T191|Tumor, Krukenberg's
C0022790|T191|Krukenbergs Tumor
C0022790|T191|Krukenberg tumor (disorder)
C1333319|T191|Ductal Breast Carcinoma with Squamous Metaplasia
C1333319|T191|Ductal Carcinoma of Breast with Squamous Metaplasia
C1333319|T191|Ductal Carcinoma of the Breast with Squamous Metaplasia
C1711312|T191|Breast Carcinoma with Osseous Metaplasia
C1335148|T191|Osteosarcoma Arising in Paget Disease of Bone
C1335148|T191|Paget's Osteosarcoma
C1335148|T191|Osteosarcoma Arising in Paget's Disease of Bone
C1335148|T191|Paget Osteosarcoma
C1335148|T191|Osteosarcoma Arising in Osteitis Deformans
C1335148|T191|Osteosarcoma Arising in Bone Paget's Disease
C1335148|T191|Osteosarcoma Arising in Osseous Paget's Disease
C1145205|T200|Zoledronic Acid
C1145205|T200|Zometa
C1145205|T200|ZOL 446
C1145205|T200|zoledronic acid
C1145205|T200|NDC-Zoledronate
C1145205|T200|Zoledronic acid
C1145205|T200|[1-Hydroxy-2-(1H-imidazol-1-yl)ethylidene]bisphosphonic Acid
C1145205|T200|ZOLEDRONIC ACID
C1145205|T200|CGP42446A
C1145205|T200|INJECTION, ZOLEDRONIC ACID (ZOMETA), 1 MG
C1145205|T200|INJECTION, ZOLEDRONIC ACID (ZOMETA), 1 MG ADMINISTERED
C1145205|T200|Reclast
C1145205|T200|CGP 42446
C1334705|T191|Metachronous Wilms Tumor
C1334705|T191|Metachronous Wilms Tumor of the Kidney
C1334705|T191|Metachronous Wilms' Tumor
CL412333|T061|Breast Irradiation
CL412333|T061|breast irradiation
C1518013|T191|Low Grade Adenosquamous Breast Carcinoma
C1518013|T191|Infiltrating Breast Syringomatous Adenoma
C100068|T061|Cardiac Ablation
C100068|T061|CATH ABLATION
C100068|T061|Catheter Ablation
C100068|T061|Ablation, Catheter
C100068|T061|Cardiac ablation
C100068|T061|ABLATION CATH
C2985560|T061|Radioembolization
C2985560|T061|intra-arterial brachytherapy
C2985560|T061|Radioembolisation
C2985560|T061|radioembolization
C2985560|T061|transarterial radioembolization
C0700596|T116|Leuprolide Acetate
C0700596|T116|D-Leu^6^, desGly-NH>2<^10^-LHRH ethylamide monoacetate
C0700596|T116|Procrin
C0700596|T116|TAP 144
C0700596|T116|Enanton
C0700596|T116|D-leu^6^, desgly-NH>2<^10^, proethylamide^9^-GnRH monoacetate
C0700596|T116|Leuprolide acetate
C0700596|T116|LEUPROLIDE ACETATE
C0700596|T116|377526
C0700596|T116|A43818
C0700596|T116|Procren
C0700596|T116|TAP144
C0700596|T116|Leuprorelin Acetate
C0700596|T116|25379
C0700596|T116|Enantone
C0700596|T116|6-D-leucine-9-(N-ethyl-L-prolinamide)-10-deglycinamide luteinizing hormone-releasing factor (pig) monoacetate
C0700596|T116|6-D-Leucine-9-(N-ethyl-L-prolinamide)-10-deglycinamide Luteinizing Hormone-Releasing Factor (Pig) Monoacetate
C0700596|T116|LEUP
C0700596|T116|Abbott-43818
C0700596|T116|Carcinil
C0700596|T116|Leuprorelin acetate (product)
C0700596|T116|Leuplin
C0700596|T116|D-Leu<sup>6</sup>, desGly-NH<sub>2</sub><sup>10</sup>-LHRH ethylamide monoacetate
C0700596|T116|Leuprolide acetate (substance)
C0700596|T116|Trenantone
C0700596|T116|Depo-Eligard
C0700596|T116|Lucrin
C0700596|T116|Viadur
C0700596|T116|Prostap
C0700596|T116|TAP-144
C0700596|T116|6-D-leucine-9-(N-ethyl-L-prolinamide)-1-9-luteinizing hormone-releasing factor (pig) monoacetate
C0700596|T116|Acetate, Leuprolide
C0700596|T116|53714-56-0
C0700596|T116|Lupron
C0700596|T116|Lupron Depot-Ped
C0700596|T116|Abbott 43818
C0700596|T116|Lupron Depot-3 Month
C0700596|T116|A 43818
C0700596|T116|leuprolide acetate
C0700596|T116|D-leu6, desgly-NH2 10, proethylamide9-GnRH monoacetate
C0700596|T116|A-43818
C0700596|T116|Leuprorelin acetate
C0700596|T116|Enantone-Gyn
C0700596|T116|Lupron Depot
C0700596|T116|Leuprolide Acetate [Chemical/Ingredient]
C0700596|T116|Lucrin Depot
C0700596|T116|D-Leu6, desGly-NH2 10-LHRH ethylamide monoacetate
C0700596|T116|Uno-Enantone
C0700596|T116|Ginecrin
C0700596|T116|74381-53-6 (acetate)
C0700596|T116|6-D-Leucine-9-(N-ethyl-L-prolinamide)-1-9-luteinizing Hormone-releasing Factor (Pig) Monoacetate
C0700596|T116|Lupron Depot-4 Month
C0700596|T116|D-leu<sup>6</sup>, desgly-NH<sub>2</sub><sup>10</sup>, proethylamide<sup>9</sup>-GnRH monoacetate
C0700596|T116|Eligard
C0861834|T191|Recurrent Malignant Duodenal Neoplasm
C0861834|T191|Malignant neoplasm of duodenum recurrent
C1336816|T191|Transplant-Related Skin Squamous Cell Carcinoma
C0743505|T190|Endocervical Mass
C0278780|T191|Recurrent Adult Acute Myeloid Leukemia
C0278780|T191|Recurrent Adult Acute Myelogenous Leukemia
C0278780|T191|relapsed adult AML
C0278780|T191|recurrent acute myeloid leukemia, adult
C0278780|T191|Relapsed Adult Acute Myelogenous Leukemia
C0278780|T191|adult acute myelogenous leukemia, relapsed
C0278780|T191|adult acute myeloid leukemia, relapsed
C0278780|T191|relapsed adult acute myelogenous leukemia
C0278780|T191|ANLL, relapsed, adult
C0278780|T191|adult acute nonlymphocytic leukemia, relapsed
C0278780|T191|myeloid leukemia, relapsed adult acute
C0278780|T191|relapsed adult ANLL
C0278780|T191|adult leukemia, relapsed acute myeloid
C0278780|T191|recurrent adult AML
C0278780|T191|AML, adult recurrent
C0278780|T191|Relapsed Adult Acute Myeloid Leukemia
C0278780|T191|recurrent adult ANLL
C0278780|T191|leukemia, relapsed adult acute nonlymphocytic
C0278780|T191|adult ANLL, recurrent
C0278780|T191|adult leukemia, relapsed acute nonlymphocytic
C0278780|T191|AML, relapsed, adult
C0278780|T191|relapsed adult acute myeloid leukemia
C0278780|T191|myelogenous leukemia, relapsed adult acute
C0278780|T191|Relapsed Adult AML
C0278780|T191|acute nonlymphocytic leukemia, relapsed, adult
C0278780|T191|recurrent adult acute myeloid leukemia
C0278780|T191|adult AML, recurrent
C0278780|T191|acute myeloid leukemia, relapsed, adult
C0278780|T191|leukemia, relapsed adult acute myeloid
C0278780|T191|acute myelogenous leukemia, relapsed, adult
C0278780|T191|Recurrent Adult Acute Non-Lymphocytic Leukemia
C0278780|T191|nonlymphocytic leukemia, relapsed adult acute
C0278780|T191|ANLL, adult recurrent
C0278780|T191|adult leukemia, relapsed acute myelogenous
C0278780|T191|leukemia, relapsed adult acute myelogenous
C0278780|T191|adult AML, relapsed
C0278780|T191|Recurrent Adult AML
C1334799|T191|Monomorphic T/NK-Cell Post-Transplant Lymphoproliferative Disorder
C1334799|T191|Monomorphic T-Cell PTLD
C1334799|T191|Monomorphic T-Cell Post-Transplant Lymphoproliferative Disorder
C0043308|T061|X-ray Therapy
C0043308|T061|x-ray therapy
C0686055|T191|Metastatic Malignant Neoplasm to the Esophagus
C0686055|T191|Metastasis to the Esophagus
C0686055|T191|Esophageal Metastasis
C0686055|T191|Metastases to the Esophagus
C0686055|T191|Metastatic Tumor to the Esophagus
C0686055|T191|Metastatic Neoplasm to the Esophagus
C0686055|T191|Metastases to Esophagus
C0686055|T191|Metastasis to Esophagus
C1334784|T191|Mixed Epithelial and Mesenchymal Hepatoblastoma
C0278553|T191|Recurrent Colon Carcinoma
C0278553|T191|Recurrent Cancer of the Colon
C0278553|T191|Colon carcinoma recurrent
C0278553|T191|Recurrent Colon Cancer
C0278553|T191|Recurrent Cancer of Colon
C0278553|T191|colon cancer, recurrent
C0278553|T191|Carcinoma colon recurrent
C0278553|T191|recurrent colon cancer
C0278553|T191|Colon cancer recurrent
C1335923|T191|Sarcomatoid Carcinoma of the Penis
C1335923|T191|Sarcomatoid Penile Squamous Cell Carcinoma
C1335923|T191|Sarcomatous Carcinoma of the Penis
C1335923|T191|Sarcomatoid Penile Carcinoma
C1335923|T191|Spindle Cell Carcinoma of the Penis
C1335923|T191|Squamous Cell Carcinoma of the Penis, Sarcomatoid Type
C1335923|T191|Squamous Cell Carcinoma of Penis, Sarcomatoid Type
C0586555|T033|Epigastric Mass
C0586555|T033|Epigastric mass (finding)
C0586555|T033|Epigastric mass
C1519358|T033|Slow Growing Mass
C1334735|T191|Metastatic Non-Cutaneous Melanoma
C0475388|T185|T2b Stage Finding
C0475388|T185|Tumour stage T2b
C0475388|T185|T2b Tumor Stage
C0475388|T185|Tumor Stage T2b
C0475388|T185|T2b Stage
C0475388|T185|T2b TNM Finding
C0475388|T185|Tumor stage T2b (finding)
C0475388|T185|T2b Primary Tumor Stage Finding
C0475388|T185|T2b Tumor Finding
C0475388|T185|T2b Primary Tumor Finding
C0475388|T185|T2b Cancer Stage Finding
C0475388|T185|T2b
C0475388|T185|Tumor stage T2b
C1541447|T191|Recurrent Childhood Grade III Lymphomatoid Granulomatosis
C0279981|T191|Childhood Fibrosarcoma
C0279981|T191|sarcoma, fibro-, childhood
C0279981|T191|fibrosarcoma, pediatric
C0279981|T191|pediatric fibrosarcoma
C0279981|T191|fibrosarcoma, childhood
C0279981|T191|Pediatric Fibrosarcoma
C0279981|T191|childhood fibrosarcoma
C0920506|T191|Environment-Related Malignant Neoplasm
C0920506|T191|Environment-Related Cancer
C0920506|T191|Environmental Malignant Neoplasm
C0920506|T191|Environmental Cancers
C0920506|T191|Environmental Cancer
C0024103|T033|Breast Lump
C0024103|T033|Unspecified lump in breast
C0024103|T033|BREAST MASS
C0024103|T033|Breast Mass
C0024103|T033|Breast lump (finding)
C0024103|T033|MASS BREAST (NOS)
C0024103|T033|area of enhancement
C0024103|T033|Breast Nodule
C0024103|T033|lesion
C0024103|T033|nodule
C0024103|T033|mass
C0024103|T033|breast mass
C0024103|T033|Lumpy breast
C0024103|T033|BREAST LUMPS
C0024103|T033|breast nodule
C0024103|T033|Breast mass NOS
C0024103|T033|Lump in Breast
C0024103|T033|Breast mass
C0024103|T033|Lumpy breasts
C0024103|T033|Mass in Breast
C0024103|T033|Breast lump NOS
C0024103|T033|breast density
C0024103|T033|Breast irregular nodularity
C0024103|T033|Breast nodule
C0024103|T033|BREAST NODULE
C0024103|T033|Lump or mass in breast
C0024103|T033|Mammary gland mass
C0024103|T033|LUMPS, BREAST
C0024103|T033|focus
C0024103|T033|nodular enhancement
C0024103|T033|Breast lump
C0024103|T033|Mass in breast
C0006098|T061|Internal Radiation Therapy
C0006098|T061|Radiation Brachytherapy
C0006098|T061|Brachytherapy, Radioisotope
C0006098|T061|Brachytherapy
C0006098|T061|BRACHYTHER RADIOISOTOPE
C0006098|T061|Contact radiation therapy procedure
C0006098|T061|Brachytherapy - action (qualifier value)
C0006098|T061|Radioisotope Brachytherapy
C0006098|T061|BRACHYTHER
C0006098|T061|Brachytherapy - action
C0006098|T061|Brachytherapy NOS
C0006098|T061|CURIETHER
C0006098|T061|Plesiotherapy radiation
C0006098|T061|Curietherapy
C0006098|T061|brachytherapy
C0006098|T061|Brachytherapy procedure
C0006098|T061|Internal Radiation Brachytherapy
C0006098|T061|radiation brachytherapy
C0006098|T061|internal radiation
C0006098|T061|Internal Radiation
C0006098|T061|RADIOISOTOPE BRACHYTHER
C0033822|T191|Pseudomyxoma Peritonei
C0033822|T191|Gelatinous Ascites
C0033822|T191|pseudomyxoma peritonei
C0033822|T191|Mucinous Ascites
C0033822|T191|Peritoneal Cavity Pseudomyxoma Peritonei
C0033822|T191|Myxoma Peritonei
C0033822|T191|Well Differentiated Peritoneal Mucinous Adenocarcinoma
C1332182|T191|Adult Anaplastic Large Cell Lymphoma
C1332182|T191|Adult CD30+ Anaplastic Large Cell Lymphoma
C1332182|T191|Adult K-1+ Anaplastic Large Cell Lymphoma
C0854746|T191|Stage III AIDS-Related Anal Canal Cancer
C0854746|T191|Stage III AIDS-Related Anal Canal Cancer AJCC v6
C0854746|T191|Stage III AIDS-Related Anal Canal Cancer AJCC v7
C1332982|T191|Childhood Mesenchymal Chondrosarcoma
C1332982|T191|Pediatric Mesenchymal Chondrosarcoma
C0278802|T191|Recurrent Uterine Corpus Carcinoma
C0278802|T191|recurrent uterine cancer
C0278802|T191|endometrial carcinoma, recurrent
C0278802|T191|carcinoma of the endometrium, recurrent
C0278802|T191|recurrent cancer of the endometrium
C0278802|T191|endometrial cancer, recurrent
C0278802|T191|Endometrial cancer recurrent
C0278802|T191|Endometrial carcinoma recurrent
C0278802|T191|recurrent carcinoma of the endometrium
C0278802|T191|cancer of the endometrium, recurrent
C0278802|T191|Carcinoma endometrial recurrent
C0278802|T191|Recurrent Endometrial Cancer
C0278802|T191|Cancer of endometrium recurrent
C0278802|T191|recurrent endometrial carcinoma
C0278802|T191|recurrent endometrial cancer
C0278802|T191|Recurrent Corpus Uteri Cancer
C0278802|T191|uterine cancer, recurrent
C0278802|T191|Recurrent Uterine Corpus Cancer
C1333006|T191|Childhood Testicular Choriocarcinoma
C1333006|T191|Pediatric Choriocarcinoma of the Testis
C1333006|T191|Childhood Choriocarcinoma of the Testis
C1333006|T191|Pediatric Choriocarcinoma of Testis
C1333006|T191|Childhood Choriocarcinoma of Testis
C1333006|T191|Pediatric Testicular Choriocarcinoma
C1332214|T191|Adult Primary Cutaneous Anaplastic Large Cell Lymphoma
C1332214|T191|Adult Primary Cutaneous CD30+ Anaplastic Large Cell Lymphoma
C1332214|T191|Adult Primary Cutaneous K-1+ Anaplastic Large Cell Lymphoma
C2985557|T061|Gamma Irradiation
C2985557|T061|gamma irradiation
C106073|T061|Double Strand Brachytherapy
C1709109|T033|N3b Stage Finding
C1709109|T033|N3b Lymph Node Stage
C1709109|T033|N3b TNM Finding
C1709109|T033|N3b
C1709109|T033|N3b Regional Lymph Node Stage Finding
C1709109|T033|N3b Node Finding
C1709109|T033|N3b Lymph Node Finding
C1709109|T033|N3b Regional Lymph Nodes Finding
C1709109|T033|Lymph Node Stage N3b
C1709109|T033|Node Stage N3b
C1709109|T033|N3b Stage
C1709109|T033|N3b Cancer Stage Finding
C1709109|T033|N3b Node Stage
C1335496|T191|Primitive Neuroectodermal Tumor with Leptomeningeal Spread
C1332967|T191|Childhood Diffuse Large B -Cell Lymphoma
C1332967|T191|Pediatric Diffuse Large B Cell Lymphoma
C1335459|T191|Postsurgical Stage II Hepatoblastoma
C1332954|T191|Childhood Central Nervous System Immature Teratoma
C115031|T191|Stage III Childhood Anaplastic Large Cell Lymphoma
C0334497|T191|Pericanalicular Fibroadenoma
C0334497|T191|Pericanalicular Fibroadenoma of the Breast
C0334497|T191|Pericanalicular Fibroadenoma of Breast
C0334497|T191|Pericanalicular fibroadenoma (morphologic abnormality)
C0334497|T191|Pericanalicular Breast Fibroadenoma
C0334497|T191|Pericanalicular fibroadenoma
C0346979|T191|Metastatic Malignant Neoplasm to the Bone Marrow
C0346979|T191|Metastatic Neoplasm to the Bone Marrow
C0346979|T191|Metastases to the Bone Marrow
C0346979|T191|Metastatic Tumor to the Bone Marrow
C0346979|T191|bone marrow metastasis
C0346979|T191|Metastasis to the Bone Marrow
C2986509|T061|Accelerated-fraction Radiation Therapy
C2986509|T061|accelerated-fraction radiation therapy
C0454077|T061|Photon Beam Radiation Therapy
C0454077|T061|Electron Beam Therapy
C0454077|T061|Teleradiotherapy using beta particles
C0454077|T061|electron beam therapy
C0454077|T061|Teleradiotherapy beta particles
C0454077|T061|photon beam radiation therapy
C0454077|T061|Teleradiotherapy using electrons (procedure)
C0454077|T061|Betatron electron teletherapy
C0454077|T061|Electron teleradiotherap
C0454077|T061|Teleradiotherapy using electrons
C0454077|T061|Electron teletherapy
C115443|T191|Recurrent Nasal Cavity and Paranasal Sinus Squamous Cell Carcinoma
CL448469|T191|Recurrent Malignant Neoplasm of Salivary Gland
C1519369|T191|Anaplastic Large Cell Lymphoma, Sarcomatoid Subtype
C0494164|T191|Metastatic Malignant Neoplasm to the Small Intestine
C0494164|T191|Secondary Malignant Neoplasm to the Small Bowel
C0494164|T191|Metastases to Small Intestine
C0494164|T191|Secondary Malignant Tumor to the Small Bowel
C0494164|T191|Secondary Malignant Tumor to the Small Intestine
C0494164|T191|Metastasis to the Small Intestine
C0494164|T191|Secondary Malignant Neoplasm to the Small Intestine
C0494164|T191|Metastatic Neoplasm to the Small Intestine
C0494164|T191|Metastasis to the Small Bowel
C1332051|T191|AIDS-Related Non-Hodgkin Lymphoma
C1332051|T191|AIDS-related NHL
C1332051|T191|AIDS-related Non-Hodgkin lymphoma
C1332051|T191|AIDS-Related Non-Hodgkin's Lymphoma
C0280386|T191|Recurrent Nasopharyngeal Keratinizing Squamous Cell Carcinoma
C0280386|T191|Relapsed Nasopharyngeal Keratinizing Epidermoid Carcinoma
C0280386|T191|Recurrent Keratinizing Epidermoid Carcinoma of Nasopharynx
C0280386|T191|Relapsed Keratinizing Epidermoid Carcinoma of Nasopharynx
C0280386|T191|nasopharynx squamous cell carcinoma, recurrent
C0280386|T191|epidermoid carcinoma of the nasopharynx, recurrent
C0280386|T191|Recurrent Keratinizing Squamous Cell Carcinoma of Nasopharynx
C0280386|T191|Relapsed Keratinizing Squamous Cell Carcinoma of the Nasopharynx
C0280386|T191|Relapsed Keratinizing Squamous Cell Carcinoma of Nasopharynx
C0280386|T191|Recurrent Nasopharyngeal Keratinizing Epidermoid Carcinoma
C0280386|T191|Relapsed Keratinizing Epidermoid Carcinoma of the Nasopharynx
C0280386|T191|Nasopharyngeal squamous cell carcinoma recurrent
C0280386|T191|Recurrent Keratinizing Epidermoid Carcinoma of the Nasopharynx
C0280386|T191|nasopharyngeal squamous cell carcinoma, recurrent
C0280386|T191|Relapsed Nasopharyngeal Keratinizing Squamous Cell Carcinoma
C0280386|T191|squamous cell carcinoma of the nasopharynx, recurrent
C0280386|T191|Recurrent Keratinizing Squamous Cell Carcinoma of the Nasopharynx
C0280386|T191|recurrent squamous cell carcinoma of the nasopharynx
C0684833|T191|Metastatic Malignant Neoplasm to the Chest Wall
C0684833|T191|Metastatic Neoplasm to the Chest Wall
C0684833|T191|Secondary Malignant Tumor to the Chest Wall
C0684833|T191|Secondary Malignant Neoplasm to the Chest Wall
C0684833|T191|Metastasis to the Chest Wall
C0684833|T191|Metastatic Tumor to the Chest Wall
C1266166|T191|Conventional Osteosarcoma
C1266166|T191|osteogenic sarcoma, undifferentiated
C1266166|T191|anaplastic osteosarcoma
C1266166|T191|Central Osteosarcoma
C1266166|T191|Central osteosarcoma (morphologic abnormality)
C1266166|T191|Intracortical Osteosarcoma
C1266166|T191|Anaplastic osteosarcoma
C1266166|T191|undifferentiated osteosarcoma
C1266166|T191|anaplastic osteogenic sarcoma
C1266166|T191|Medullary osteosarcoma
C1266166|T191|osteosarcoma, undifferentiated
C1266166|T191|intracortical osteosarcoma
C1266166|T191|Central osteosarcoma
C1266166|T191|Intracortical Osteogenic Sarcoma
C1266166|T191|Conventional Central Osteosarcoma
C1266166|T191|sarcoma, osteogenic anaplastic
C1266166|T191|sarcoma, osteogenic undifferentiated
C1266166|T191|undifferentiated osteogenic sarcoma
C1266166|T191|central osteosarcoma
C1266166|T191|Intracortical osteosarcoma (morphologic abnormality)
C1266166|T191|osteosarcoma, anaplastic
C1266166|T191|Intracortical osteosarcoma
C1266166|T191|Medullary Osteosarcoma
C1266166|T191|osteogenic sarcoma, anaplastic
C1266166|T191|Conventional central osteosarcoma
C0398434|T060|Axillary Lymph Node Biopsy
C0398434|T060|Axillary Node Biopsy
C0398434|T060|axillary node biopsy
C0398434|T060|axillary lymph node biopsy
C0398434|T060|Biopsy of axillary lymph node (procedure)
C0398434|T060|Biopsy of axillary lymph node
C1332288|T191|Secondary Supratentorial Anaplastic Astrocytoma
C1332288|T191|Anaplastic Secondary Supratentorial Astrocytoma
C1332288|T191|Grade III Secondary Supratentorial Astrocytic Tumor
C1332288|T191|Grade III Secondary Supratentorial Astrocytoma
C1332288|T191|Undifferentiated Secondary Supratentorial Astrocytoma
C1332288|T191|Grade III Secondary Supratentorial Astrocytic Neoplasm
C115206|T033|Cognitive Side Effects of Cancer Therapy
C0278696|T191|Stage I Childhood Hepatocellular Carcinoma
C0278696|T191|Stage I Childhood Hepatocellular Carcinoma AJCC v7
C0278696|T191|Stage I Childhood Hepatocellular Carcinoma AJCC v6
C0278696|T191|Stage I Childhood Hepatoma
C0278696|T191|Stage I Pediatric Liver Cell Carcinoma
C0278696|T191|stage I childhood liver cancer
C0278696|T191|Stage I Childhood Liver Cell Carcinoma
C0278696|T191|Stage I Pediatric Hepatocellular Carcinoma
C0278696|T191|Stage I Pediatric Hepatoma
C1335519|T191|Acinar Prostate Adenocarcinoma, Sarcomatoid Variant
C1335519|T191|Sarcomatoid Carcinoma of the Prostate
C1335519|T191|Prostate Carcinosarcoma
C1335519|T191|Sarcomatoid Carcinoma of Prostate
C1335519|T191|Prostate Sarcomatoid Carcinoma
C115357|T191|Recurrent Childhood Anaplastic Large Cell Lymphoma
C115357|T191|recurrent childhood anaplastic large cell lymphoma
C0494165|T191|Metastatic Malignant Neoplasm to the Liver
C0494165|T191|Liver Metastases
C0494165|T191|Metastatic Tumor to the Liver
C0494165|T191|Metastatic Neoplasm to the Liver
C0494165|T191|Metastases to liver, NOS
C0494165|T191|liver metastasis
C0494165|T191|Liver Metastasis
CL447336|T061|Mesh Brachytherapy
C1879503|T061|AC Regimen
C1879503|T061|Adriamycin-Cytoxan Regimen
C1879503|T061|CA Regimen
C1879503|T061|AC regimen
C1879503|T061|AC
C1879503|T061|Adriamycin-cyclophosphamide regimen
C1334685|T191|Medulloblastoma with Leptomeningeal Spread
C1514835|T191|Renal Cell Carcinoma with Constitutional Chromosome 3 Translocations
C3272623|T201|Deep Adventitial Inked Margin
C1709263|T191|Nonestrogen-Dependent Cancer
C1709263|T191|Nonestrogen-Dependent Carcinoma
C1517029|T033|Extensive Necrosis
C1301090|T201|Size of base of tumor at cut edge, after sectioning
C1301090|T201|Size of base of tumor at cut edge, after sectioning (observable entity)
C1301090|T201|Size of base of tumour at cut edge, after sectioning
C0259785|T191|Anaplastic (Malignant) Meningioma
C0259785|T191|Malignant Meningioma
C0259785|T191|MENINGIOMA, ANAPLASTIC, MALIGNANT
C0259785|T191|malignant meningioma
C0259785|T191|ANAPLASTIC MENINGIOMA
C0259785|T191|Anaplastic Meningioma
C0259785|T191|MENINGIOMA, MALIGNANT
C0259785|T191|Meningioma, Malignant
C0259785|T191|MALIGNANT MENINGIOMA
CL448449|T191|Recurrent Extranodal Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue
CL448449|T191|Recurrent Extranodal Marginal Zone B-Cell Lymphoma (MALT Type)
CL448449|T191|Relapsed Extranodal Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue
CL448449|T191|Recurrent Extranodal Marginal Zone B-Cell Lymphoma of Mucosa-Associated Lymphoid Tissue
CL448449|T191|Relapsed MALT Type Extranodal Marginal Zone B-Cell Lymphoma
C0334500|T191|Giant Fibroadenoma
C0334500|T191|Giant Fibroadenoma of the Breast
C0334500|T191|Giant fibroadenoma (morphologic abnormality)
C0334500|T191|[M]Giant fibroadenoma
C0334500|T191|Serocystic disease of Brodie
C0334500|T191|Giant fibroadenoma
C0334500|T191|[M] Giant fibroadenoma
C0334500|T191|Giant fibroadenoma of breast
C0334500|T191|Giant Fibroadenoma of Breast
C0334500|T191|Giant fibroadenoma of breast (disorder)
C1707604|T049|Cytosine to Adenosine Transversion Abnormality
C1707604|T049|Cytosine to Adenosine Transversion
C1707604|T049|Cytosine to Adenosine Mutation
C1334990|T033|Non-Metastatic Mass
C1334990|T033|Nonmetastatic Mass
C114759|T191|Childhood Brain Stem Gliosarcoma
C114759|T191|gliosarcoma, childhood brain stem
C114759|T191|childhood brain stem gliosarcoma
C114759|T191|childhood brainstem gliosarcoma
C114759|T191|gliosarcoma, childhood brainstem
C1710406|T049|Thymidine to Guanosine Transversion Abnormality
C1710406|T049|Thymidine to Guanosine Transversion
C1710406|T049|Thymidine to Guanosine Mutation
C0279602|T191|Fibroblastic Osteosarcoma
C0279602|T191|fibroblastic osteosarcoma
C0279602|T191|osteosarcoma, fibrosarcomatous
C0279602|T191|sarcoma, osteogenic fibroblastic
C0279602|T191|fibrosarcomatous osteosarcoma
C0279602|T191|Fibroblastic osteosarcoma
C0279602|T191|Fibrosarcomatous Osteosarcoma
C0279602|T191|Osteofibrosarcoma
C0279602|T191|Fibrosarcomatous Osteogenic Sarcoma
C0279602|T191|fibrosarcomatous osteogenic sarcoma
C0279602|T191|osteosarcoma, fibroblastic
C0279602|T191|osteogenic sarcoma, fibrosarcomatous
C0279602|T191|Fibroblastic osteosarcoma (morphologic abnormality)
C0279602|T191|fibroblastic osteogenic sarcoma
C0279602|T191|osteogenic sarcoma, fibroblastic
C0279602|T191|Fibroblastic Osteogenic Sarcoma
C0278586|T191|Metastatic Ewing Sarcoma
C0278586|T191|metastatic tumors of the Ewing's family
C0278586|T191|metastatic Ewing's sarcoma
C0278586|T191|Ewing's tumour metastatic
C0278586|T191|Ewing's sarcoma metastatic
C0278586|T191|Ewing's sarcoma, metastatic
C0278586|T191|Ewing's Sarcoma, Metastatic
C0278586|T191|Metastatic Ewing's Sarcoma
C0278586|T191|Ewing's tumor metastatic
C1518574|T191|Oncocytic Breast Carcinoma
CL412338|T061|Partial Breast Irradiation
CL412338|T061|partial breast irradiation
C1963256|T046|Ulceration
C1963256|T046|Ulceration Adverse Event
C1963256|T046|Ulcus
C1963256|T046|Ulcer
C1963256|T046|Ulcerative lesion
C1963256|T046|Ulceration (qualifier value)
C1963256|T046|ulcer
C1963256|T046|Ulcer [Disease/Finding]
C1963256|T046|Ulcer NOS
C1963256|T046|Ulcerated
C1963256|T046|Ulcers
C1963256|T046|Ulcerative (qualifier value)
C1963256|T046|Ulcer (morphologic abnormality)
C1963256|T046|Ulcer (disorder)
C1963256|T046|ulceration
C1963256|T046|Ulcerative
C1963256|T046|Ulcer - lesion
C1963256|T046|ULCER
C1963256|T046|ULCERATION
C1963256|T046|Ulcerating
C1334036|T191|Hodgkin-Like Post-Transplant Lymphoproliferative Disorder
C1334036|T191|Hodgkin lymphoma-like post-transplant lymphoproliferative disorder
C1334036|T191|Hodgkin's-Like Post-Transplant Lymphoproliferative Disorder
C1334036|T191|Hodgkin-like PTLD
C1334036|T191|Hodgkin lymphoma - like PTLD
C1334036|T191|Hodgkin's-like PTLD
C0205697|T191|Sarcomatoid Carcinoma
C0205697|T191|spindle cell squamous carcinoma
C0205697|T191|Sarcomatoid carcinoma
C0205697|T191|PSEUDOSARCOMATOUS CARCINOMA
C0205697|T191|SPINDLE CELL CARCINOMA
C0205697|T191|Carcinomas, Spindle-Cell
C0205697|T191|Spindle cell carcinoma
C0205697|T191|Spindle cell carcinoma (morphologic abnormality)
C0205697|T191|sarcomatoid carcinoma
C0205697|T191|Spindle-Cell Carcinomas
C0205697|T191|Spindle-Cell Carcinoma
C0205697|T191|CARCINOMA, SPINDLE CELL, MALIGNANT
C0205697|T191|Pseudosarcoma
C0205697|T191|Spindle Cell Carcinoma
C0205697|T191|Spindle cell carcinoma, NOS
C0205697|T191|Pseudosarcomatous carcinoma (morphologic abnormality)
C0205697|T191|polypoid carcinoma
C0205697|T191|Carcinoma, Spindle Cell
C0205697|T191|Carcinoma, Spindle-Cell
C0205697|T191|pseudosarcoma
C0205697|T191|Pseudosarcomatous Carcinoma
C0205697|T191|Pseudosarcomatous carcinoma
C0205697|T191|spindle cell carcinoma
C0281642|T191|Childhood Acute Myeloid Leukemia with Minimal Differentiation
C0281642|T191|Childhood Acute Myeloid Leukemia Minimally Differentiated
C0281642|T191|M0 Childhood Acute Minimally Differentiated Myeloid Leukemia
C0281642|T191|Childhood Acute Minimally Differentiated Myeloid Leukemia (M0)
C0281642|T191|M0 Pediatric Acute Minimally Differentiated Myeloid Leukemia
C0281642|T191|Pediatric Acute Minimally Differentiated Myeloid Leukemia
C0281642|T191|Pediatric Acute M0 Leukemia
C0281642|T191|Childhood Acute M0 Leukemia
C0281642|T191|Childhood Acute Minimally Differentiated Myeloid Leukemia
CL412303|T061|Pretargeted Radioimmunotherapy
CL412303|T061|pretargeted radioimmunotherapy
C1334750|T191|Methotrexate-Associated Peripheral T-Cell Lymphoma
C0008994|T121|Clodronate Disodium
C0008994|T121|CL2MDP
C0008994|T121|Clodronate disodium (product)
C0008994|T121|Clasteon
C0008994|T121|disodium dichloromethylene diphosphonate
C0008994|T121|Disodium, Clodronate
C0008994|T121|clodronate disodium
C0008994|T121|Clodronate disodium (substance)
C0008994|T121|Sodium, Clodronate
C0008994|T121|Clodronate Sodium
C0008994|T121|Ossiten
C0008994|T121|Dichloromethylene Diphosphonate
C0008994|T121|Bonefos
C0008994|T121|Sodium clodronate
C0008994|T121|CLODRONATE DISODIUM
C0008994|T121|clodronic acid, disodium salt
C0008994|T121|clodronate
C0008994|T121|Clodronate (substance)
C0008994|T121|Loron
C0008994|T121|Mebonat
C0008994|T121|Disodium clodronate
C0008994|T121|Clodronate
C0008994|T121|Clodronic Acid Disodium Salt
C0008994|T121|713466
C0008994|T121|Difosfonal
C0008994|T121|Clodronate disodium
C1709094|T049|Multiple Transversion Abnormalities
C1709094|T049|Multiple Transversion Mutations
C1709094|T049|Transversion Mutations
C0001632|T061|Adrenalectomy
C0001632|T061|Excision of adrenal gland
C0001632|T061|Adrenalectomy (procedure)
C0001632|T061|Adrenalectomies
C0001632|T061|ADRENALECTOMY
C0001632|T061|Adrenal Gland Excision
C0001632|T061|Adrenalectomy NOS
C0001632|T061|Excision of Adrenal Gland
C0001632|T061|Excision of adrenal gland operations
C0001632|T061|adrenalectomy
C1332977|T191|Childhood Leukemia
C1332977|T191|Leukemia, Childhood
C0342500|T047|Adrenal Mass
C0342500|T047|Adrenal mass
C0342500|T047|Mass of adrenal gland
C0342500|T047|Mass of adrenal gland (finding)
C1541316|T191|Adult Giant Cell Glioblastoma
C1541316|T191|giant cell glioblastoma, adult
C1541316|T191|adult giant cell glioblastoma
C1336024|T191|Solar Radiation-Related Skin Squamous Cell Carcinoma
C1335505|T191|Prostate Carcinoma Metastatic to the Bone
C0475393|T185|Tumor stage T3bii
C0475393|T185|Tumour stage T3bii
C0475393|T185|Tumor stage T3bii (finding)
C1335721|T191|Recurrent Urinary Tract Carcinoma
C1335721|T191|Recurrent Urinary Tract Cancer
C0475398|T185|T4d Stage Finding
C0475398|T185|T4d Cancer Stage Finding
C0475398|T185|T4d Stage
C0475398|T185|T4d Tumor Stage
C0475398|T185|Tumour stage T4d
C0475398|T185|T4d Tumor Finding
C0475398|T185|Tumor Stage T4d
C0475398|T185|T4d Primary Tumor Finding
C0475398|T185|T4d Primary Tumor Stage Finding
C0475398|T185|T4d TNM Finding
C0475398|T185|Tumor stage T4d (finding)
C0475398|T185|T4d
C0475398|T185|Tumor stage T4d
C0445306|T082|Wart size
C0445306|T082|Wart size (observable entity)
C0445306|T082|Size of warts
C1334740|T191|Metastatic Signet Ring Cell Breast Carcinoma
C1334740|T191|Metastatic Mammary Signet Ring Cell Carcinoma
C1334740|T191|Metastatic Signet Ring Cell Carcinoma of Breast
C1334740|T191|Metastatic SRC Carcinoma of Breast
C1334740|T191|Metastatic SRC Carcinoma of the Breast
C1334740|T191|Metastatic Signet Ring Cell Carcinoma of the Breast
C1334740|T191|Metastatic SRC Breast Carcinoma
C0684550|T191|Metastatic Malignant Neoplasm to the Spine
C0684550|T191|Metastatic Cancer to the Spine
C0684550|T191|Metastasis to the Spine
C0684550|T191|Metastatic Tumor to the Vertebral Column
C0684550|T191|Metastatic Neoplasm to the Spine
C0684550|T191|Metastasis to Spine
C0684550|T191|Metastases to Spine
C0684550|T191|Metastatic Neoplasm to the Vertebral Column
C0684550|T191|Metastases to the Spine
C0684550|T191|Metastatic Cancer to the Vertebral Column
C0684550|T191|Metastatic Tumor to the Spine
C0677964|T046|Unresectable Mass
C0854858|T191|Recurrent T Lymphoblastic Leukemia/Lymphoma
C0854858|T191|Relapsed Precursor T Lymphoblastic Lymphoma/Leukemia
C0854858|T191|Recurrent Precursor T-Lymphoblastic Lymphoma/Leukemia
C0117339|T121|Toremifene Citrate
C0117339|T121|FC 1157a
C0117339|T121|FC-1157a
C0117339|T121|FC1157a
C0117339|T121|toremifene citrate
C0117339|T121|Fareston
C0117339|T121|2-(p-[(Z)-4-chloro-1,2-diphenyl-1-butenyl]-phenoxy)- N,N-dimethylethylamine citrate (1:1)
C0117339|T121|TOREMIFENE CITRATE
C0117339|T121|Acapodene
C0117339|T121|(Z)-2-[4-(4-Chloro-1,2-diphenyl-1-butenyl)phenoxy]-N,N-dimethylethanamine 2-Hydroxy-1,2,3-propanetricarboxylate (1:1)
C0117339|T121|Toremifene Citrate [Chemical/Ingredient]
C0117339|T121|Toremifene citrate (product)
C0117339|T121|Toremifene citrate (substance)
C0117339|T121|Toremifene citrate
C0117339|T121|GTx-006
C0117339|T121|Citrate, Toremifene
C0117339|T121|Toremifene Citrate (1:1)
C1334813|T191|Mucoepidermoid Breast Carcinoma
C1334813|T191|Mucoepidermoid Carcinoma of the Breast
C1334813|T191|Mucoepidermoid Carcinoma of Breast
C0862435|T191|Recurrent Renal Cell Carcinoma
C0862435|T191|Renal carcinoma recurrent
C0862435|T191|recurrent hypernephroma
C0862435|T191|hypernephroma, recurrent
C0862435|T191|Carcinoma kidney recurrent
C0862435|T191|Kidney cancer recurrent
C0862435|T191|Kidney carcinoma recurrent
C0862435|T191|recurrent renal cell carcinoma
C0862435|T191|Renal cancer recurrent
C0862435|T191|kidney cancer, recurrent
C0862435|T191|Renal Cell Carcinoma, Recurrent
C0862435|T191|renal cell cancer, recurrent
C0862435|T191|Hypernephroma recurrent
C0862435|T191|Renal cell carcinoma recurrent
C0862435|T191|recurrent kidney cancer
C0862435|T191|recurrent renal cell cancer
C0862435|T191|Relapsed Renal Cell Carcinoma
C0862435|T191|renal cell carcinoma, recurrent
C0281706|T191|Stage IV Childhood Burkitt Lymphoma
C0281706|T191|Stage IV Childhood Burkitt's Lymphoma
C0281706|T191|Stage IV Pediatric Small Non-Cleaved Cell Lymphoma
C0281706|T191|Metastatic Pediatric Small Non-Cleaved Cell Lymphoma
C0281706|T191|Pediatric Small Non-Cleaved Cell Lymphoma Stage IV
C0281706|T191|Stage IV Childhood Small Non-Cleaved Cell Lymphoma
C0281706|T191|Childhood Small Non-Cleaved Cell Lymphoma Stage IV
C0281706|T191|Metastatic Childhood Small Non-Cleaved Cell Lymphoma
C0023488|T191|Radiation-Related Leukemia
C0023488|T191|Radiation-Induced Leukemia
C0746319|T033|Positive Lymph Node
C0746319|T033|node-positive
C0854849|T191|Recurrent Mycosis Fungoides
C0854849|T191|Relapsed Mycosis Fungoides
C0854849|T191|Mycosis fungoides recurrent
C0854849|T191|Mycosis Fungoides Recurrent
C0854849|T191|Mycosis Fungoides Relapsed
C0015133|T121|Etoposide
C0015133|T121|ETOPOSIDE
C0015133|T121|VP-16-213
C0015133|T121|4'-Demethylepipodophyllotoxin 9-[4,6-O-ethylidene-beta-D-glucopyranoside]
C0015133|T121|Vepesid
C0015133|T121|VP-16
C0015133|T121|EPEG
C0015133|T121|Toposar
C0015133|T121|etoposide
C0015133|T121|Lastet
C0015133|T121|Demethyl Epipodophyllotoxin Ethylidine Glucoside
C0015133|T121|9-[(4,6-O-Ethylidene-beta-D-glucopyranosyl]oxy)-5,8,8a,9-tetrahydro-5-(4-hydroxy-3,5-dimethoxyphenyl)furo[3',4':6,7]naphtho[2,3-d]-1,3-dioxol-6(5aH)-one
C0015133|T121|VP 16-213
C0278785|T191|Recurrent Adult Acute Lymphoblastic Leukemia
C0278785|T191|acute lymphocytic leukemia, recurrent, adult
C0278785|T191|Relapsed Adult Acute Lymphoblastic Leukemia
C0278785|T191|recurrent adult ALL
C0278785|T191|leukemia, relapsed adult acute lymphocytic
C0278785|T191|relapsed adult ALL
C0278785|T191|lymphocytic leukemia, relapsed adult acute
C0278785|T191|Relapsed Adult Acute Lymphogenous Leukemia
C0278785|T191|ALL, relapsed, adult
C0278785|T191|Recurrent Adult Precursor Lymphoblastic Leukemia
C0278785|T191|Relapsed Adult Acute Lymphoid Leukemia
C0278785|T191|acute lymphocytic leukemia, relapsed, adult
C0278785|T191|relapsed ALL, adult
C0278785|T191|Recurrent Adult Acute Lymphocytic Leukemia
C0278785|T191|ALL, recurrent, adult
C0278785|T191|recurrent adult acute lymphocytic leukemia
C0278785|T191|recurrent ALL, adult
C0278785|T191|recurrent adult acute lymphoblastic leukemia
C0278785|T191|adult acute lymphocytic leukemia, relapsed
C0278785|T191|Recurrent Adult Acute Lymphoid Leukemia
C0278785|T191|Relapsed Adult ALL
C0278785|T191|Relapsed Adult Acute Lymphocytic Leukemia
C0278785|T191|relapsed adult acute lymphocytic leukemia
C0278785|T191|Recurrent Adult ALL
C0278785|T191|Recurrent Adult Acute Lymphogenous Leukemia
CL454080|T191|Glioblastoma by Gene Expression Profile
C2985435|T049|Founder Mutation
C2985435|T049|founder mutation
C1334441|T191|Lung Carcinoma Metastatic to the Brain
C1519485|T191|Squamous Cell Breast Carcinoma, Acantholytic Variant
C1510796|T191|Adenosquamous Breast Carcinoma
C116445|T061|Computed Tomography-Guided Optical Sensor-Guided Radiofrequency Ablation
C0278737|T191|Stage III Childhood Lymphoblastic Lymphoma
C0278737|T191|Childhood Lymphoblastic Lymphoma Stage III
C0278737|T191|Pediatric Lymphoblastic Lymphoma Stage III
C0278737|T191|Stage III Childhood Precursor Lymphoblastic Lymphoma
C0278737|T191|Stage III Pediatric Lymphoblastic Lymphoma
C0685120|T191|Metastatic Malignant Neoplasm to the Pericardium
C0685120|T191|Metastatic Neoplasm to the Pericardium
C0001688|T169|Side Effect
C0001688|T169|undesirable effects
C0001688|T169|side effect
C0001688|T169|Treatment Side Effects
C0001688|T169|injurious effects
C0001688|T169|ADV EFF
C0001688|T169|adverse effects
C0001688|T169|side effects
C0001688|T169|AE
C0854920|T191|Recurrent Ureter Carcinoma
C0854920|T191|Ureter cancer recurrent
C0854920|T191|Relapsed Ureter Cancer
C0854920|T191|Relapsed Cancer of the Ureter
C0854920|T191|Recurrent Ureter Cancer
C0854920|T191|Ureteric Cancer, Recurrent
C0854920|T191|Malignant neoplasm of ureter recurrent
C0854920|T191|Relapsed Ureteral Cancer
C0854920|T191|Relapsed Cancer of Ureter
C0854920|T191|Ureteric cancer recurrent
CL055234|T191|Recurrent Ewing Sarcoma/Peripheral Primitive Neuroectodermal Tumor
CL055234|T191|Recurrent Tumors of Ewing's Family
CL055234|T191|Recurrent Tumors of the Ewing's Family
CL055234|T191|Recurrent Ewing's Sarcoma/Peripheral Primitive Neuroectodermal Tumor
C0280376|T191|Recurrent Oropharyngeal Squamous Cell Carcinoma
C0280376|T191|Recurrent Oropharyngeal Epidermoid Carcinoma
C0280376|T191|Relapsed Squamous Cell Carcinoma of Oropharynx
C0280376|T191|Recurrent Oropharyngeal SCC
C0280376|T191|Recurrent Epidermoid Carcinoma of Oropharynx
C0280376|T191|Recurrent Squamous Cell Carcinoma of Oropharynx
C0280376|T191|Relapsed SCC of the Oropharynx
C0280376|T191|epidermoid carcinoma of the oropharynx, recurrent
C0280376|T191|squamous cell carcinoma of the oropharynx, recurrent
C0280376|T191|Relapsed Oropharyngeal Squamous Cell Carcinoma
C0280376|T191|Oropharyngeal squamous cell carcinoma recurrent
C0280376|T191|Recurrent SCC of the Oropharynx
C0280376|T191|Relapsed Epidermoid Carcinoma of the Oropharynx
C0280376|T191|oropharyngeal squamous cell carcinoma, recurrent
C0280376|T191|Recurrent Squamous Cell Carcinoma of the Oropharynx
C0280376|T191|Relapsed Squamous Cell Carcinoma of the Oropharynx
C0280376|T191|Relapsed SCC of Oropharynx
C0280376|T191|Recurrent SCC of Oropharynx
C0280376|T191|oropharynx squamous cell carcinoma, recurrent
C0280376|T191|Relapsed Oropharyngeal SCC
C0280376|T191|Recurrent Epidermoid Carcinoma of the Oropharynx
C0280376|T191|recurrent squamous cell carcinoma of the oropharynx
C0280376|T191|Relapsed Epidermoid Carcinoma of Oropharynx
C0280376|T191|Relapsed Oropharyngeal Epidermoid Carcinoma
C0445034|T033|M0 Stage Finding
C0445034|T033|M0 TNM Finding
C0445034|T033|M0 category (finding)
C0445034|T033|Metastasis Stage M0
C0445034|T033|M0 Distant Metastasis Finding
C0445034|T033|M0 category
C0445034|T033|M0 distant metastasis stage
C0445034|T033|M0 Cancer Stage Finding
C0445034|T033|M0 Metastasis Stage
C0445034|T033|M0 Metastasis Finding
C0445034|T033|Metastasis stage M0
C0445034|T033|M0 Distant Metastasis Stage Finding
C0445034|T033|M0 Stage
C0445034|T033|M0
C0445034|T033|M0 stage
C1516823|T049|Embryonic Lethal Mutation
C1516823|T049|Embryonic Lethal Mutation Abnormality
CL472853|T191|Refractory Childhood Hodgkin Lymphoma
C0280098|T191|Undifferentiated Carcinoma of Unknown Primary
C1519478|T049|Splice-Site Mutation
C1519478|T049|Intron Splice Site Mutation
C1519478|T049|Splice-Site Mutation Abnormality
C1519478|T049|Splice-Juction Mutation
C1519478|T049|Intronic Splice Site Mutation
C0886487|T191|Recurrent Childhood Malignant Germ Cell Neoplasm
C0886487|T191|recurrent childhood malignant germ cell tumor
C0886487|T191|germ cell tumor, recurrent, childhood
C0886487|T191|recurrent germ cell tumor, childhood
C0886487|T191|recurrent childhood germ cell tumor
C0886487|T191|Recurrent Childhood Malignant Germ Cell Tumor
C0886487|T191|pediatric recurrent germ cell tumor
C0886487|T191|recurrent germ cell tumor, pediatric
C0886487|T191|germ cell tumor, recurrent, pediatric
C1711276|T191|Lung Carcinosarcoma
C0280734|T191|AIDS-Related Malignant Neoplasm
C0280734|T191|AIDS-Related Malignancy
C0280734|T191|AIDS Related Cancer
C0280734|T191|AIDS-Related Cancer
C0280734|T191|AIDS-Related Malignancies
C0280734|T191|AIDS-related cancer
C2985434|T049|Disease-causing Mutation
C2985434|T049|disease-causing mutation
C1336922|T191|AIDS-Related Burkitt Lymphoma with Plasmacytoid Differentiation
C1336922|T191|AIDS-Related Burkitt's Lymphoma with Plasmacytoid Differentiation
C1511281|T191|Breast Adenocarcinoma with Spindle Cell Metaplasia
CL421682|T061|Palliative Radiation Therapy
CL421682|T061|palliative radiation therapy
C1334440|T191|Lung Carcinoma Metastatic to the Bone
C1831915|T061|Hyperfractionation
C1831915|T061|Hyperfractionated Radiation Therapy
C1831915|T061|superfractionated radiation therapy
C1831915|T061|hyperfractionated radiation therapy
C1831915|T061|hyperfractionation
C1831915|T061|Hyperfractionated Radiation
C1527223|T121|Paclitaxel Albumin-Stabilized Nanoparticle Formulation
C1527223|T121|protein-bound paclitaxel
C1527223|T121|Abraxane
C1527223|T121|Nanoparticle Albumin-bound Paclitaxel
C1527223|T121|Albumin-bound Paclitaxel
C1527223|T121|nab-paclitaxel
C1527223|T121|ABI-007
C1527223|T121|Nanoparticle Paclitaxel
C1527223|T121|Albumin-Stabilized Nanoparticle Paclitaxel
C1527223|T121|paclitaxel albumin-stabilized nanoparticle formulation
C1527223|T121|ABI 007
C1527223|T121|nanoparticle paclitaxel
C0860594|T191|Metastatic Melanoma
C0860594|T191|Malignant melanoma, metastatic
C0860594|T191|Metastatic malignant melanoma (disorder)
C0860594|T191|Metastatic malignant melanoma
C0860594|T191|melanoma, metastatic
C0860594|T191|Malignant melanoma, metastatic (morphologic abnormality)
C0860594|T191|metastatic melanoma
C0860594|T191|Metastatic melanoma
C1334736|T191|Metastatic Ovarian Small Cell Carcinoma, Hypercalcemic Type
CL472835|T191|Recurrent Pancreatic Neuroendocrine Carcinoma
C0153687|T191|Metastatic Malignant Neoplasm to the Skin
C0153687|T191|Metastases to Skin
C0153687|T191|Metastases to skin, NOS
C0153687|T191|Skin Metastasis
C0153687|T191|Metastatic Tumor to the Skin
C0153687|T191|Metastasis to Skin
C0153687|T191|Skin Metastases
C0153687|T191|Metastatic Neoplasm to the Skin
C1334277|T191|Invasive Ductal and Lobular Carcinoma
C1334277|T191|Infiltrating Ductal and Lobular Carcinoma
C1334277|T191|Invasive Duct and Lobular Carcinoma
C0278746|T191|Recurrent Vaginal Carcinoma
C0278746|T191|Recurrent Vagina Cancer
C0278746|T191|Relapsed Vagina Cancer
C0278746|T191|Recurrent Cancer of the Vagina
C0278746|T191|Recurrent Cancer of Vagina
C0278746|T191|Relapsed Cancer of Vagina
C0278746|T191|vagina cancer, recurrent
C0278746|T191|Vaginal cancer recurrent
C0278746|T191|recurrent carcinoma of the vagina
C0278746|T191|Relapsed Vaginal Cancer
C0278746|T191|vaginal cancer, recurrent
C0278746|T191|Relapsed Cancer of the Vagina
C0278746|T191|Cancer of vagina recurrent
C0278746|T191|cancer of the vagina, recurrent
C0278746|T191|Recurrent Vaginal Cancer
C0278746|T191|recurrent cancer of the vagina
C0278746|T191|recurrent vaginal cancer
C0278746|T191|carcinoma of the vagina, recurrent
C0278746|T191|recurrent vagina cancer
CL433902|T191|Recurrent Childhood Anaplastic Astrocytoma
CL433902|T191|recurrent childhood anaplastic astrocytoma
C0677779|T191|Hereditary Wilms Tumor
C0677779|T191|Familiar Wilms Tumor
C0677779|T191|Familial Wilms' Tumor
C0677779|T191|Familial Wilms Tumor
C0677779|T191|Wilms tumor, familial
C0677779|T191|Hereditary Nephroblastoma (WT1)
C0677779|T191|hereditary Wilms' tumor (WT1)
C0677779|T191|Hereditary Renal Adenosarcoma (WT1)
C0677779|T191|hereditary Wilms tumor
C0677779|T191|Hereditary Kidney Adenosarcoma (WT1)
C0677779|T191|Hereditary Wilms' Tumor (WT1)
C0677779|T191|Hereditary Wilms' Tumor
C0861212|T191|Recurrent Centroblastic Lymphoma
C0861212|T191|Centroblastic lymphoma recurrent
C0577731|T191|Disseminated Adenocarcinoma
C0577731|T191|Disseminated adenocarcinoma (morphologic abnormality)
C0577731|T191|Disseminated adenocarcinoma
C2986685|T191|Stage III AIDS-Related Lymphoma
C2986685|T191|stage III AIDS-related lymphoma
C1370446|T191|Recurrent Plasma Cell Myeloma
C1370446|T191|Recurrent Multiple Myeloma
C1370446|T191|Plasma cell myeloma recurrent
C1332972|T191|Childhood Infratentorial Ependymoblastoma
C1332972|T191|Pediatric Infratentorial Ependymoblastoma
C1442161|T045|Gene Deletion
C1442161|T045|Gene Deletions
C1442161|T045|Gene deletion
C1442161|T045|gene deletion mutation
C1442161|T045|Gene deletion (attribute)
C1442161|T045|Deletion
C1442161|T045|MOLPATH.DEL
C1442161|T045|Deletion, Gene
C1442161|T045|gene deletion
C1442161|T045|Deletions, Gene
C1442161|T045|Gene Deletion Abnormality
C0441961|T033|N3 Stage Finding
C0441961|T033|N3 Node Finding
C0441961|T033|N3 Regional Lymph Node Stage Finding
C0441961|T033|N3 lymph node stage
C0441961|T033|N3 Node Stage
C0441961|T033|N3 Cancer Stage Finding
C0441961|T033|Node Stage N3
C0441961|T033|N3 Lymph Node Stage
C0441961|T033|N3 stage
C0441961|T033|N3 TNM Finding
C0441961|T033|N3 category
C0441961|T033|Node stage N3
C0441961|T033|N3 category (finding)
C0441961|T033|N3
C0441961|T033|N3 Stage
C0441961|T033|Lymph Node Stage N3
C0441961|T033|N3 Regional Lymph Nodes Finding
C0441961|T033|N3 Lymph Node Finding
C3272450|T033|N1bIII Stage Finding
C0346997|T191|Metastatic Malignant Neoplasm to the Vagina
C0346997|T191|Metastatic Neoplasm to the Vagina
C0346997|T191|Metastasis to the Vagina
C0346997|T191|Secondary Tumor to Vagina
C0346997|T191|Metastasis to Vagina
C0346997|T191|Secondary Tumor to the Vagina
C0677898|T191|Invasive Malignant Neoplasm
C0677898|T191|Infiltrating Malignant Neoplasm
C0677898|T191|invasive cancer
C0677898|T191|infiltrating cancer
C0030185|T191|Paget Disease of the Breast
C0030185|T191|Paget's Disease of the Breast
C0030185|T191|Mammary Paget's Disease
C0030185|T191|Paget's Disease of Breast
C1333988|T191|Hereditary Male Breast Carcinoma
C1333988|T191|Familial Male Breast Carcinoma
C2919520|T081|Calculated volume of neoplasm based on largest dimension using magnetic resonance imaging
C2919520|T081|Calculated volume of neoplasm based on largest dimension using magnetic resonance imaging (observable entity)
C1332270|T191|Paget Disease of the Anal Margin
C1332270|T191|Perianal Skin Paget's Disease
C1332270|T191|Paget's Disease of the Anal Margin
C1332270|T191|Anal Margin Paget's Disease
C1300943|T201|Tumor size, non-dominant nodule, greatest dimension
C1300943|T201|Tumor size, non-dominant nodule, greatest dimension (observable entity)
C1300943|T201|Tumour size, non-dominant nodule, greatest dimension
C0206629|T191|Pulmonary Blastoma
C0206629|T191|Blastomas, Pulmonary
C0206629|T191|pulmonary blastoma
C0206629|T191|PULM BLASTOMAS
C0206629|T191|Blastoma of the Lung
C0206629|T191|BLASTOMA PULM
C0206629|T191|PULM BLASTOMA
C0206629|T191|BLASTOMAS PULM
C0206629|T191|Blastoma of Lung
C0206629|T191|Pulmonary blastoma
C0206629|T191|Pneumoblastoma
C0206629|T191|Pulmonary Blastomas
C0206629|T191|Pulmonary blastoma (morphologic abnormality)
C0206629|T191|Lung Blastoma
C0206629|T191|[M] Pulmonary blastoma
C0206629|T191|[M]Pulmonary blastoma
C0206629|T191|Pulmonary Blastoma [Disease/Finding]
C0206629|T191|Blastoma, Pulmonary
C2919402|T033|Largest dimension of in situ neoplasm
C2919402|T033|Largest dimension of in situ neoplasm (observable entity)
C1368019|T191|Paget Disease
C1368019|T191|Paget's Cell Neoplasm
C1368019|T191|Paget disease
C1368019|T191|Paget's Disease
C1368019|T191|Paget Cell Neoplasm
C1960177|T191|Colonic Mass
C1960177|T191|Colonic mass
C1960177|T191|Neoplasm of colon
C1960177|T191|Neoplasm of the Colon
C1960177|T191|Neoplasm, Colon
C1960177|T191|Mass of colon (finding)
C1960177|T191|colon neoplasm
C1960177|T191|Tumor of Colon
C1960177|T191|Neoplasm of colon (disorder)
C1960177|T191|colon tumor or cancer
C1960177|T191|Colon Tumor
C1960177|T191|COLONIC NEOPLASM
C1960177|T191|Neoplasms, Colon
C1960177|T191|Neoplasm of Colon
C1960177|T191|Colonic Tumor
C1960177|T191|COLON TUMOR
C1960177|T191|Colonic Neoplasms
C1960177|T191|NEOPL COLONIC
C1960177|T191|Colon neoplasm
C1960177|T191|Neoplasm, Colonic
C1960177|T191|Colonic Neoplasm
C1960177|T191|Tumor of colon
C1960177|T191|Tumour of colon
C1960177|T191|Colonic neoplasm NOS
C1960177|T191|NEOPLASM OF COLON
C1960177|T191|Tumor of the Colon
C1960177|T191|Mass of colon
C1960177|T191|COLONIC NEOPL
C1960177|T191|Neoplasms, Colonic
C1960177|T191|Colon neoplasm NOS
C1960177|T191|Colon neoplasia
C1960177|T191|Colonic tumor
C1960177|T191|Colon Neoplasm
C1960177|T191|Colon Neoplasms
C1960177|T191|COLON NEOPL
C1960177|T191|Colonic Neoplasms [Disease/Finding]
C1333137|T191|Complex Fibroadenoma
C1333137|T191|Complex Fibroadenoma of the Breast
C1333137|T191|Complex Fibroadenoma of Breast
C115381|T191|Recurrent Childhood Supratentorial Primitive Neuroectodermal Tumor
C115381|T191|recurrent neuroblastoma, pediatric cerebral
C115381|T191|recurrent pediatric supratentorial PNET
C115381|T191|recurrent primitive neuroectodermal tumor, pediatric supratentorial
C115381|T191|pediatric supratentorial primitive neuroectodermal tumor, recurrent
C115381|T191|recurrent neuroblastoma, childhood cerebral
C115381|T191|recurrent pediatric cerebral neuroblastoma
C115381|T191|PNET, recurrent childhood supratentorial
C115381|T191|recurrent neuroectodermal tumor, pediatric, primitive, supratentorial
C115381|T191|childhood supratentorial primitive neuroectodermal tumor, recurrent
C115381|T191|pediatric cerebral neuroblastoma, recurrent
C115381|T191|recurrent primitive neuroectodermal tumor, supratentorial, pediatric
C115381|T191|recurrent PNET, childhood supratentorial
C115381|T191|recurrent childhood supratentorial primitive neuroectodermal tumor
C115381|T191|recurrent supratentorial primitive neuroectodermal tumor, childhood
C115381|T191|PNET, recurrent pediatric supratentorial
C115381|T191|recurrent childhood supratentorial primitive neuroectodermal tumors
C115381|T191|cerebral neuroblastoma, recurrent, childhood
C115381|T191|recurrent primitive neuroectodermal tumor, childhood supratentorial
C115381|T191|recurrent cerebral neuroblastoma, pediatric
C115381|T191|recurrent neuroblastoma, cerebral, pediatric
C115381|T191|childhood cerebral neuroblastoma, recurrent
C115381|T191|cerebral neuroblastoma, recurrent, pediatric
C115381|T191|recurrent childhood cerebral neuroblastoma
C115381|T191|pediatric supratentorial PNET, recurrent
C115381|T191|recurrent neuroblastoma, cerebral, childhood
C115381|T191|recurrent cerebral neuroblastoma, childhood
C115381|T191|childhood supratentorial PNET, recurrent
C115381|T191|recurrent pediatric supratentorial primitive neuroectodermal tumors
C115381|T191|recurrent pediatric primitive neuroectodermal tumor, supratentorial
C115381|T191|recurrent PNET, pediatric supratentorial
C115381|T191|recurrent pediatric supratentorial primitive neuroectodermal tumor
C115381|T191|recurrent supratentorial primitive neuroectodermal tumor, pediatric
C115381|T191|PNET, supratentorial, childhood, recurrent
C115381|T191|recurrent neuroectodermal tumor, childhood, primitive, supratentorial
C115381|T191|recurrent childhood supratentorial PNET
C115381|T191|recurrent primitive neuroectodermal tumor, supratentorial, childhood
C115381|T191|PNET, supratentorial, pediatric, recurrent
C115381|T191|recurrent childhood primitive neuroectodermal tumor, supratentorial
C1519218|T191|Secondary Prostate Urothelial Carcinoma
C0278870|T191|Recurrent Uveal Melanoma
C0278870|T191|uveal melanoma, recurrent
C0278870|T191|recurrent uveal melanoma
C0278870|T191|recurrent intraocular melanoma
C0278870|T191|Recurrent Melanoma of Uvea
C0278870|T191|Recurrent Melanoma of the Uvea
C0278870|T191|intraocular melanoma, recurrent
C0278870|T191|melanoma, uveal recurrent
C1710108|T033|Slow Growing Painless Mass
C0279917|T191|Stage IV Childhood Hodgkin Lymphoma
C0279917|T191|Pediatric Hodgkin's Disease Stage IV
C0279917|T191|stage IV childhood Hodgkin lymphoma
C0279917|T191|Pediatric Hodgkin's Lymphoma Stage IV
C0279917|T191|Stage IV Childhood Hodgkin's Lymphoma
C0279917|T191|Childhood Hodgkin's Lymphoma Stage IV
C0279917|T191|Stage IV Pediatric Hodgkin Lymphoma
C0279917|T191|Childhood Hodgkin's Disease Stage IV
C0279917|T191|Stage IV Pediatric Hodgkin's Lymphoma
C3282903|T191|Metastatic Carcinoma to the Liver
C1879758|T191|Atypical Medullary Breast Carcinoma
C1879758|T191|Infiltrating Ductal Breast Carcinoma with Medullary Features
C0054427|T061|CAF Regimen
C0054427|T061|Cyclophosphamide-Adriamycin-Fluorouracil regimen
C0054427|T061|CAF regimen
C0054427|T061|CAFFI
C0054427|T061|FAC protocol
C0054427|T061|CDF
C0054427|T061|Cyclophosphamide/Doxorubicin/Fluorouracil
C0054427|T061|CAF protocol
C0054427|T061|FAC
C0054427|T061|CAF
C0054427|T061|CTX/DOX/5-FU
C0054427|T061|Cyclophosphamide-Adriamycin-Fluorouracil Regimen
C1709611|T191|Radiation-Related Osteosarcoma
C1709611|T191|Postradiation Osteosarcoma
C1514169|T191|Pleomorphic Breast Carcinoma
C1514169|T191|Anaplastic Breast Carcinoma
C1518010|T061|Low Dose Radiation Therapy
C1518010|T061|Low Dose Radiation
C1332966|T191|Childhood Desmoplastic Small Round Cell Tumor
C1332966|T191|Pediatric Desmoplastic Small Round Cell Tumor
C1332966|T191|small round cell tumor, desmoplastic, childhood
C1332966|T191|Desmoplastic Small Round-Cell Tumor
C1332966|T191|childhood desmoplastic small round cell tumor
C1332966|T191|tumor, desmoplastic small round cell, childhood
C1332966|T191|DSRCT
C1332966|T191|Desmoplastic Small Round Cell Tumor
C1332966|T191|Desmoplastic Small Round-Cell Neoplasm
C1511760|T045|Deletion Mutation
C1511760|T045|deletion
C1511760|T045|Deletion Abnormality
C1511760|T045|Deletion
C1511760|T045|Mutations, Deletion
C1511760|T045|Deletion Mutations
C1511760|T045|Mutation, Deletion
C0345960|T191|Lung Giant Cell Carcinoma
C0345960|T191|Giant Cell Carcinoma of Lung
C0345960|T191|Giant cell carcinoma of lung (disorder)
C0345960|T191|Giant cell carcinoma of lung
C0345960|T191|Giant Cell Carcinoma of the Lung
C1334280|T191|Invasive Papillary Breast Carcinoma
C1334280|T191|Invasive papillary breast carcinoma
C1334280|T191|Infiltrating Papillary Breast Carcinoma
C1334746|T191|Methotrexate-Associated Diffuse Large B-Cell Lymphoma
CL388411|T061|Accelerated Radiation Therapy
CL388411|T061|accelerated radiation therapy
CL374463|T061|Laser Interstitial Thermal Therapy
CL374463|T061|laser interstitial thermal therapy
CL374463|T061|LITT
CL454081|T191|Proneural Glioblastoma
C0085203|T061|Radiosurgery
C0085203|T061|Stereo radiosurgery NOS
C0085203|T061|stereotaxic radiation therapy
C0085203|T061|STEREOTACTIC RADIOSURG
C0085203|T061|Stereotactic radiosurgery (procedure)
C0085203|T061|Stereotactic Radiotherapy
C0085203|T061|SBRT
C0085203|T061|Radiosurgeries
C0085203|T061|Stereotactic External Beam Irradiation
C0085203|T061|Radiosurgery, Stereotactic
C0085203|T061|RADIOSURG STEREOTACTIC
C0085203|T061|stereotaxic radiosurgery
C0085203|T061|Stereotactic radiosurgery, not otherwise specified
C0085203|T061|Stereotactic Radiation Therapy
C0085203|T061|Stereotactic Radiosurgery
C0085203|T061|radiosurgery
C0085203|T061|stereotactic body radiation therapy
C0085203|T061|RADIOSURG
C0085203|T061|Radiation Surgery
C0085203|T061|Stereotactic radiosurgery
C0085203|T061|Radiosurgeries, Stereotactic
C0085203|T061|radiation surgery
C0085203|T061|Stereotactic Radiosurgeries
C0085203|T061|stereotactic radiation therapy
C0085203|T061|stereotactic external-beam radiation therapy
C0085203|T061|stereotactic radiosurgery
C0236022|T191|Aggravated Malignant Neoplasm
C0236022|T191|Malignant neoplasm aggravated
C0236022|T191|Neoplasm malignant aggravated
C0278738|T191|Stage IV Childhood Lymphoblastic Lymphoma
C0278738|T191|Metastatic Childhood Lymphoblastic Lymphoma
C0278738|T191|Childhood Stage IV Lymphoblastic Lymphoma
C0278738|T191|Stage IV Pediatric Lymphoblastic Lymphoma
C0278738|T191|Stage IV Childhood Precursor Lymphoblastic Lymphoma
C0278738|T191|Metastatic Pediatric Lymphoblastic Lymphoma
C0278738|T191|Childhood Lymphoblastic Lymphoma Stage IV
C0278738|T191|Pediatric Lymphoblastic Lymphoma Stage IV
C0278738|T191|Pediatric Stage IV Lymphoblastic Lymphoma
C0279634|T191|Childhood Acute Myeloid Leukemia without Maturation
C0279634|T191|Pediatric AML without Maturation
C0279634|T191|M1 Childhood Acute Myeloid Leukemia without Maturation
C0279634|T191|Childhood Acute Myelocytic Leukemia without Maturation
C0279634|T191|M1 Childhood Acute Myelocytic Leukemia without Maturation
C0279634|T191|M1 childhood acute myeloblastic leukemia without maturation
C0279634|T191|Childhood Acute Myelogenous Leukemia without Maturation
C0279634|T191|childhood AML without maturation
C0279634|T191|Childhood Acute M1 Leukemia
C0279634|T191|pediatric acute myeloblastic leukemia without maturation
C0279634|T191|M1 childhood AML without maturation
C0279634|T191|Pediatric Acute Myeloblastic Leukemia without Maturation
C0279634|T191|Childhood Acute Myeloblastic Leukemia without Maturation
C0279634|T191|M1 Pediatric Acute Myelogenous Leukemia without Maturation
C0279634|T191|M1 pediatric acute myeloblastic leukemia without maturation
C0279634|T191|childhood acute M1 leukemia
C0279634|T191|Pediatric Acute Myelogenous Leukemia without Maturation
C0279634|T191|M1 Childhood Acute Myelogenous Leukemia without Maturation
C0279634|T191|M1 Pediatric Acute Myelocytic Leukemia without Maturation
C0279634|T191|M1 Pediatric Acute Myeloblastic Leukemia without Maturation
C0279634|T191|Pediatric Acute Myelocytic Leukemia without Maturation
C0279634|T191|childhood acute myeloblastic leukemia without maturation (M1)
C0279634|T191|Childhood Acute Myeloblastic Leukemia Without Maturation (M1)
C0279634|T191|Pediatric Acute Myeloid Leukemia without Maturation
C0279634|T191|M1 leukemia, childhood acute
C0279634|T191|M1 Pediatric Acute Myeloid Leukemia without Maturation
C0279634|T191|pediatric acute M1 leukemia
C0279634|T191|Childhood AML without Maturation
C0279634|T191|M1 Pediatric Acute Myelogenous Leukemia
C0279634|T191|M1 Childhood Acute Myeloblastic Leukemia without Maturation
C0279634|T191|Pediatric Acute M1 Leukemia
C0546540|T061|Right Radical Mastectomy
C494392|T116|Denosumab
C494392|T116|AMG-162
C494392|T116|Denosumab (product)
C494392|T116|Xgeva
C494392|T116|Densosumab
C494392|T116|Prolia
C494392|T116|DENOSUMAB
C494392|T116|denosumab
C494392|T116|Denosumab (substance)
C494392|T116|AMG 162
C0862636|T191|Metastatic Prostatic Adenocarcinoma
C0862636|T191|Adenocarcinoma of the prostate metastatic
CL448424|T191|Recurrent Melanoma of the Skin
CL448424|T191|Recurrent Malignant Skin Melanoma
CL448424|T191|Recurrent Cutaneous Melanoma
CL448424|T191|Recurrent Melanoma of Skin
CL448424|T191|Recurrent Malignant Melanoma of the Skin
CL448424|T191|Recurrent Malignant Melanoma of Skin
C2986677|T191|Stage I Childhood Non-Hodgkin Lymphoma
C2986677|T191|stage I childhood non-Hodgkin lymphoma
C0804677|T081|Tumor Size
C0804677|T081|tumor size
C0804677|T081|Tumor size
C0804677|T081|Size:Len:Pt:Tumor:Qn
C0804677|T081|Tumor size (observable entity)
C0804677|T081|Size Tumor
C0804677|T081|size of tumor
C0804677|T081|Size:Length:Point in time:Tumor:Quantitative
C0804677|T081|Tumour size
C0804677|T081|Size of tumor
C0804677|T081|Size of tumour
C1321870|T191|Childhood Extraocular Retinoblastoma
C1321870|T191|pediatric extraocular retinoblastoma
C1321870|T191|childhood extraocular retinoblastoma
C1321870|T191|Pediatric Extraocular Retinoblastoma
C3273255|T049|Unmutated Immunoglobulin Heavy Chain Variable Region Gene
C1300453|T201|Tumor size, dominant nodule
C1300453|T201|Tumor size, dominant nodule (observable entity)
C1300453|T201|Tumour size, dominant nodule
C0861555|T191|Recurrent Malignant Oral Neoplasm
C0861555|T191|Oral neoplasm malignant recurrent
C0546541|T061|Left Radical Mastectomy
C0862967|T191|Recurrent Cholangiocarcinoma
C0862967|T191|Cholangiocarcinoma recurrent
C0862967|T191|Recurrent Cholangiocellular Carcinoma
C0086330|T074|Gamma Knife
C0086330|T074|Gamma Radiosurgical Stereotactic Systems
C0086330|T074|Gamma Systems
C0086330|T074|GAMMA KNIFE RADIOSURG
C0086330|T074|Stereotactic Systems, Radiosurgical, Gamma
C0086330|T074|RADIOSURG GAMMA KNIFE
C0086330|T074|Radiosurgery, Gamma Knife
C0086330|T074|Radiosurgical Units, Stereotactic, Gamma
C0086330|T074|Gamma Knife Radiosurgery
C0086330|T074|Radiosurgeries, Gamma Knife
C0086330|T074|Gamma Knife Radiosurgeries
C0086330|T074|Stereotactic Radiosurgical Systems, Gamma
C0086330|T074|Stereotactic Systems, Frame-Guided, Radiosurgical, Gamma
C0086330|T074|Gamma Knife (physical object)
C0086330|T074|Radiosurgery using Gamma irradiation
C0086330|T074|Gamma Knives
C0086330|T074|Gamma Knife therapy
C0086330|T074|Gamma Frame-Guided Radiosurgical Stereotactic Systems
C0086330|T074|Gamma Radiosurgical Systems, Stereotactic
C1334718|T191|Metastatic Ewing Sarcoma/Peripheral Primitive Neuroectodermal Tumor
C1334718|T191|Metastatic Ewing's Sarcoma/Peripheral Primitive Neuroectodermal Tumor
C0441971|T033|Metastasis stage M1
C0441971|T033|M1 Stage Finding
C0441971|T033|M1 Distant Metastasis Stage Finding
C0441971|T033|Metastasis Stage M1
C0441971|T033|M1
C0441971|T033|M1 Metastasis Finding
C0441971|T033|M1 Metastasis Stage
C0441971|T033|M1 category
C0441971|T033|M1 category (finding)
C0441971|T033|M1 distant metastasis stage
C0441971|T033|M1 Distant Metastasis Finding
C0441971|T033|M1 Cancer Stage Finding
C0441971|T033|M1 stage
C0441971|T033|M1 Stage
C0441971|T033|M1 TNM Finding
C0278827|T191|Recurrent Bladder Carcinoma
C0278827|T191|recurrent bladder cancer
C0278827|T191|Bladder carcinoma recurrent
C0278827|T191|Relapsed Cancer of Urinary Bladder
C0278827|T191|Recurrent Bladder Cancer
C0278827|T191|Relapsed Urinary Bladder Cancer
C0278827|T191|Relapsed Cancer of the Urinary Bladder
C0278827|T191|bladder cancer, recurrent
C0278827|T191|Relapsed Bladder Cancer
C0278827|T191|Recurrent Urinary Bladder Cancer
C0278827|T191|Bladder Carcinoma Recurrent
C0278827|T191|recurrent carcinoma of the bladder
C0278827|T191|Recurrent Cancer of the Urinary Bladder
C0278827|T191|cancer of the bladder, recurrent
C0278827|T191|Relapsed Cancer of Bladder
C0278827|T191|carcinoma of the bladder, recurrent
C0278827|T191|Recurrent Cancer of Urinary Bladder
C0278827|T191|Bladder cancer recurrent
C0278827|T191|Relapsed Cancer of the Bladder
C0278827|T191|Carcinoma bladder recurrent
C0278827|T191|Recurrent Cancer of the Bladder
C0278827|T191|Urinary bladder carcinoma recurrent
C0278827|T191|Bladder Cancer, Recurrent
C0278827|T191|Carcinoma urinary bladder recurrent
C0278827|T191|recurrent cancer of the bladder
C0278827|T191|Recurrent Cancer of Bladder
C1333838|T191|Grade 2 Invasive Breast Carcinoma
C1333838|T191|Intermediate Combined Histologic Grade Infiltrating Breast Carcinoma
C1333838|T191|Moderately Differentiated Infiltrating Breast Carcinoma
C1333838|T191|Moderately Differentiated Invasive Breast Carcinoma
C1333838|T191|Grade 2 Infiltrating Breast Carcinoma
C1333838|T191|Moderately Favorable Infiltrating Breast Carcinoma
C1321722|T191|Acute Myeloid Leukemia Arising from Previous Myelodysplastic Syndrome
C1321722|T191|Acute Myeloid Leukemia with Multilineage Dysplasia following Myelodysplastic Syndrome
C1321722|T191|AML/MDS
C0948715|T033|Infusion-Related Reaction
C0948715|T033|Infusion Related Reaction
C0948715|T033|Infusion related reaction
CL448388|T191|Paget Disease of the Scrotum
CL448388|T191|Paget's Disease of Scrotum
CL448388|T191|Scrotal Paget's Disease
CL448388|T191|Paget's Disease of the Scrotum
C1332674|T191|AIDS-Related Anal Non-Hodgkin Lymphoma
C1332674|T191|AIDS-Related Anal Non-Hodgkin's Lymphoma
C1332674|T191|AIDS-Related Primary Anal Non-Hodgkin's Lymphoma
C0445039|T033|Metastasis stage MX
C0445039|T033|Metastasis Stage MX
C0445039|T033|MX Stage Finding
C0445039|T033|MX Distant Metastasis Finding
C0445039|T033|MX TNM Finding
C0445039|T033|MX Metastasis Finding
C0445039|T033|MX category
C0445039|T033|MX
C0445039|T033|MX distant metastasis stage
C0445039|T033|MX Cancer Stage Finding
C0445039|T033|MX Distant Metastasis Stage Finding
C0445039|T033|MX Stage
C0445039|T033|MX Metastasis Stage
C0445039|T033|MX category (finding)
C0445039|T033|MX stage
C1704328|T191|Osteoblastic Osteosarcoma
C1704328|T191|sarcoma, osteogenic osteoblastic
C1704328|T191|Osteoblastic sarcoma
C1704328|T191|osteogenic sarcoma, osteoblastic
C1704328|T191|Osteoblastic osteosarcoma
C1704328|T191|osteoblastic osteogenic sarcoma
C1704328|T191|osteoblastic osteosarcoma
C1704328|T191|osteosarcoma, osteoblastic
C1302656|T201|Primary tumor size
C1302656|T201|Primary tumor size (observable entity)
C1302656|T201|Primary tumour size
CL107025|T191|Metastatic Malignant Neoplasm
CL107025|T191|metastatic cancer
CL107025|T191|cancer, metastatic
CL107025|T191|Metastatic Cancer
CL107025|T191|Metastatic cancer
C2985551|T061|Charged-particle Radiation Therapy
C2985551|T061|charged-particle radiation therapy
C0445081|T033|N2c Stage Finding
C0445081|T033|N2c Node Stage
C0445081|T033|Lymph Node Stage N2c
C0445081|T033|N2c Cancer Stage Finding
C0445081|T033|N2c Lymph Node Finding
C0445081|T033|Node stage N2c (finding)
C0445081|T033|N2c Regional Lymph Nodes Finding
C0445081|T033|N2c Stage
C0445081|T033|N2c Node Finding
C0445081|T033|N2c Regional Lymph Node Stage Finding
C0445081|T033|Node Stage N2c
C0445081|T033|N2c
C0445081|T033|Node stage N2c
C0445081|T033|N2c Lymph Node Stage
C0445081|T033|N2c TNM Finding
C1333309|T191|Distantly Metastatic Malignant Neoplasm
CL433913|T191|Recurrent Childhood Glioblastoma
CL433913|T191|recurrent childhood glioblastoma
C1708261|T049|Guanosine to Adenosine Transition Abnormality
C1708261|T049|Guanosine to Adenosine Mutation
C1708261|T049|Guanosine to Adenosine Transition
C0743497|T047|Endobronchial Mass
C0079083|T197|Carboplatin
C0079083|T197|Carboplatin Hexal
C0079083|T197|Novoplatinum
C0079083|T197|Blastocarb
C0079083|T197|Carbosol
C0079083|T197|Carbosin
C0079083|T197|(SP-4-2)-diammine[1,1-cyclobutanedicarboxylato(2--)-O,O']platinum
C0079083|T197|Nealorin
C0079083|T197|cis-diammine(cyclobutanedicarboxylato)platinum II
C0079083|T197|CBDCA
C0079083|T197|1,1-cyclobutanedicarboxylic acid platinum complex
C0079083|T197|Displata
C0079083|T197|Ercar
C0079083|T197|Paraplatin
C0079083|T197|Paraplatine
C0079083|T197|platinum, diammine(1,1-cyclobutanedicarboxylato(2-))-, (SP-4-2)
C0079083|T197|Carboplatino
C0079083|T197|Paraplat
C0079083|T197|Paraplatin AQ
C0079083|T197|Carboplat
C0079083|T197|Cis-Diammine(cyclobutane-1,1-dicarboxylato)platinum
C0079083|T197|Carbotec
C0079083|T197|Platinwas
C0079083|T197|JM-8
C0079083|T197|Ribocarbo
C0079083|T197|carboplatin
C0079083|T197|CARBOPLATIN
C0079083|T197|cis-diammine(1,1-cyclobutanedicarboxylato) platinum(II)
C3274709|T191|Contralateral Breast Carcinoma
C0684572|T191|Metastatic Malignant Neoplasm to the Sternum
C0684572|T191|Metastatic Neoplasm to the Sternum
C0684572|T191|Metastatic Malignant Tumor to the Sternum
C0684572|T191|Metastasis to the Sternum
C0684572|T191|Metastatic Tumor to the Sternum
C1707256|T033|Cancer TNM Vessel Invasion Finding Category
C0671970|T114|Capecitabine
C0671970|T114|capecitabine
C0671970|T114|Xeloda
C0671970|T114|Capecitabine (substance)
C0671970|T114|capecitabine [Chemical/Ingredient]
C0671970|T114|Capecitabine (product)
C0671970|T114|5'-Deoxy-5-fluoro-N-[(pentyloxy)carbonyl]-cytidine
C0671970|T114|Ro 09-1978/000
C0671970|T114|712807
C0671970|T114|CAPECITABINE
C0671970|T114|N(4)-pentyloxycarbonyl-5'-deoxy-5-fluorocytidine
C0671970|T114|154361-50-9
C0671970|T114|CAPE
C1511305|T191|Breast Columnar Cell Mucinous Carcinoma
C0279818|T191|Recurrent Laryngeal Carcinoma
C0279818|T191|Relapsed Carcinoma of Larynx
C0279818|T191|Recurrent Carcinoma of the Larynx
C0279818|T191|Relapsed Laryngeal Carcinoma
C0279818|T191|Larynx neoplasm malignant recurrent
C0279818|T191|Laryngeal cancer recurrent
C0279818|T191|Recurrent Larynx Cancer
C0279818|T191|Recurrent Larynx Carcinoma
C0279818|T191|larynx cancer, recurrent
C0279818|T191|Relapsed Carcinoma of the Larynx
C0279818|T191|laryngeal cancer, recurrent
C0279818|T191|Relapsed Larynx Carcinoma
C0279818|T191|Malignant neoplasm of larynx recurrent
C0279818|T191|recurrent laryngeal cancer
C0279818|T191|Recurrent Carcinoma of Larynx
C0279818|T191|Recurrent Laryngeal Cancer
C0279818|T191|Larynx cancer recurrent
C0278697|T191|Stage II Childhood Hepatocellular Carcinoma
C0278697|T191|Stage II Pediatric Hepatocellular Carcinoma
C0278697|T191|Stage II Childhood Hepatoma
C0278697|T191|Stage II Pediatric Hepatoma
C0278697|T191|stage II childhood liver cancer
C0278697|T191|Stage II Childhood Liver Cell Carcinoma
C0278697|T191|Stage II Childhood Hepatocellular Carcinoma AJCC v6
C0278697|T191|Stage II Childhood Hepatocellular Carcinoma AJCC v7
C0278697|T191|Stage II Pediatric Liver Cell Carcinoma
C1112459|T191|Non-Resectable Hepatocellular Carcinoma
C490728|T121|Lapatinib
C490728|T121|GW-572016
C490728|T121|GSK572016
C490728|T121|N-(3-chloro-4-(((3-fluorobenzyl)oxy)phenyl)-6-(5-(((2-methylsulfonyl)ethyl)amino)methyl) -2-furyl)-4-quinazolinamine
C490728|T121|lapatinib
C490728|T121|GW 2016
C490728|T121|Lapatinib (substance)
C490728|T121|Lapatinib (product)
C490728|T121|GW572016
C490728|T121|LAPATINIB
C490728|T121|GW2016
C490728|T121|lapatinib [Chemical/Ingredient]
C490728|T121|GW 572016
C1711397|T191|Lung Pleomorphic Carcinoma
CL446010|T061|Scanning Proton Beam Therapy
C1334703|T191|Metachronous Malignant Neoplasm
C1334411|T191|Locally Metastatic Malignant Neoplasm
C1334411|T191|regional cancer
C2986678|T191|Stage II Childhood Non-Hodgkin Lymphoma
C2986678|T191|stage II childhood non-Hodgkin lymphoma
C562840|T191|Hereditary Breast Carcinoma
C562840|T191|Familial cancer of breast
C562840|T191|Familial cancer of breast (disorder)
C562840|T191|Familial Cancer of Breast
C562840|T191|BREAST CANCER, FAMILIAL
C562840|T191|Familial Breast Carcinoma
C562840|T191|Familial Cancer of the Breast
C562840|T191|Breast Cancer, Familial
C562840|T191|Hereditary Breast Cancer
C104933|T061|Volume Modulated Arc Therapy
C104933|T061|VMAT
C1709051|T049|Mixed Nucleotide Abnormalities
C1709051|T049|Mixed Mutations
C1709051|T049|Mixed Nucleotide Mutations
C1332990|T191|Childhood Ovarian Immature Teratoma
C1332990|T191|Pediatric Ovarian Immature Teratoma
C1332990|T191|Childhood Immature Teratoma of the Ovary
C1332990|T191|Pediatric Immature Teratoma of the Ovary
C1332990|T191|Childhood Immature Teratoma of Ovary
C1332990|T191|Pediatric Immature Teratoma of Ovary
C0338342|T191|Recurrent Childhood Medulloblastoma
C0338342|T191|PNET, infratentorial, childhood, recurrent
C0338342|T191|PNET, pediatric infratentorial, recurrent
C0338342|T191|recurrent cerebellar PNET, pediatric
C0338342|T191|recurrent cerebellar, pediatric, PNET
C0338342|T191|recurrent cerebellar PNET, childhood
C0338342|T191|recurrent cerebellar, childhood, PNET
C0338342|T191|recurrent medulloblastoma, pediatric
C0338342|T191|PNET, childhood infratentorial, recurrent
C0338342|T191|recurrent primitive neuroectodermal tumor, pediatric cerebellar
C0338342|T191|recurrent pediatric cerebellar primitive neuroectodermal tumor
C0338342|T191|recurrent PNET, pediatric infratentorial
C0338342|T191|recurrent PNET, infratentorial, pediatric
C0338342|T191|pediatric medulloblastoma, recurrent
C0338342|T191|recurrent PNET, childhood cerebellar
C0338342|T191|recurrent PNET, childhood infratentorial
C0338342|T191|recurrent medulloblastoma, childhood
C0338342|T191|recurrent PNET, infratentorial, childhood
C0338342|T191|Relapsed Pediatric Medulloblastoma
C0338342|T191|recurrent primitive neuroectodermal tumor, childhood cerebellar
C0338342|T191|childhood cerebellar PNET, recurrent
C0338342|T191|recurrent infratentorial primitive neuroectodermal tumor, childhood
C0338342|T191|pediatric infratentorial PNET, recurrent
C0338342|T191|recurrent pediatric cerebellar PNET
C0338342|T191|medulloblastoma, childhood, recurrent
C0338342|T191|recurrent infratentorial primitive neuroectodermal tumor, pediatric
C0338342|T191|childhood infratentorial primitive neuroectodermal tumor, recurrent
C0338342|T191|Relapsed Childhood Medulloblastoma
C0338342|T191|recurrent childhood medulloblastoma
C0338342|T191|recurrent childhood cerebellar PNET
C0338342|T191|recurrent pediatric infratentorial primitive neuroectodermal tumor
C0338342|T191|recurrent cerebellar primitive neuroectodermal tumor, pediatric
C0338342|T191|PNET, infratentorial, pediatric, recurrent
C0338342|T191|recurrent childhood cerebellar primitive neuroectodermal tumor
C0338342|T191|recurrent pediatric medulloblastoma
C0338342|T191|PNET, pediatric cerebellar, recurrent
C0338342|T191|childhood medulloblastoma, recurrent
C0338342|T191|childhood infratentorial PNET, recurrent
C0338342|T191|Recurrent Pediatric Medulloblastoma
C0338342|T191|recurrent cerebellar primitive neuroectodermal tumor, childhood
C0338342|T191|recurrent primitive neuroectodermal tumor, pediatric infratentorial
C0338342|T191|medulloblastoma, pediatric, recurrent
C0338342|T191|recurrent infratentorial PNET, pediatric
C0338342|T191|recurrent infratentorial, pediatric, PNET
C0338342|T191|PNET, childhood cerebellar, recurrent
C0338342|T191|PNET, cerebellar, pediatric, recurrent
C0338342|T191|recurrent infratentorial, childhood, PNET
C0338342|T191|recurrent primitive neuroectodermal tumor, childhood infratentorial
C0338342|T191|recurrent childhood infratentorial PNET
C0338342|T191|pediatric cerebellar PNET, recurrent
C0338342|T191|PNET, cerebellar, childhood, recurrent
C0338342|T191|recurrent pediatric infratentorial PNET
C0338342|T191|recurrent PNET, pediatric cerebellar
C0338342|T191|recurrent infratentorial PNET, childhood
C0338342|T191|recurrent childhood infratentorial primitive neuroectodermal tumor
C3275044|T061|Ablation of Cardiac Atrioventricular Node
C3275044|T061|ABLATION, AV NODE
C1880405|T061|Doxorubicin-Docetaxel Regimen
C1880405|T061|Adriamycin-Taxotere Regimen
C0278695|T191|Recurrent Neuroblastoma
C0278695|T191|Neuroblastoma recurrent
C0278695|T191|Relapsed Neuroblastoma
C0278695|T191|neuroblastoma, recurrent
C0278695|T191|recurrent neuroblastoma
C1332837|T191|Cancer with Regional Lymph Node Involvement
C0855078|T191|Recurrent Mixed Cellularity Classical Hodgkin Lymphoma
C0855078|T191|Relapsed Mixed Cellularity Hodgkin's Disease
C0855078|T191|Hodgkin's disease mixed cellularity recurrent
C0855078|T191|Recurrent Mixed Cellularity Hodgkin Lymphoma
C0855078|T191|Relapsed Mixed Cellularity Hodgkin's Lymphoma
C0855078|T191|Recurrent Mixed Cellularity Hodgkin's Lymphoma
C0855078|T191|Recurrent Mixed Cellularity Hodgkin's Disease
C3272440|T033|N0 (i-) Stage Finding
C2986682|T191|Locally Recurrent Malignant Neoplasm
C2986682|T191|Locally Recurrent Cancer
C2986682|T191|locally recurrent cancer
C0184913|T061|Re-Excision
C0184913|T061|Reexcision
C0686402|T191|Metastatic Malignant Neoplasm to the Brain Stem
C0686402|T191|Metastatic Neoplasm to the Brain Stem
C0686402|T191|Metastatic Tumor to the Brain Stem
C0686402|T191|Metastatic Tumor to the Brainstem
C0686402|T191|Metastatic Neoplasm to the Brainstem
C0855174|T191|Recurrent Bladder Adenocarcinoma
C0855174|T191|Relapsed Adenocarcinoma of Urinary Bladder
C0855174|T191|Bladder Adenocarcinoma, Recurrent
C0855174|T191|Recurrent Urinary Bladder Adenocarcinoma
C0855174|T191|Recurrent Adenocarcinoma of Bladder
C0855174|T191|Relapsed Adenocarcinoma of the Bladder
C0855174|T191|Relapsed Urinary Bladder Adenocarcinoma
C0855174|T191|Relapsed Adenocarcinoma of the Urinary Bladder
C0855174|T191|Recurrent Adenocarcinoma of the Bladder
C0855174|T191|Recurrent Adenocarcinoma of Urinary Bladder
C0855174|T191|Recurrent Adenocarcinoma of the Urinary Bladder
C0855174|T191|Relapsed Bladder Adenocarcinoma
C0855174|T191|Bladder adenocarcinoma recurrent
C0855174|T191|Relapsed Adenocarcinoma of Bladder
CL374485|T191|Childhood B Acute Lymphoblastic Leukemia with t(9;22)(q34;q11.2); BCR-ABL1
CL374485|T191|Childhood B-Cell Acute Lymphoblastic Leukemia with t(9;22)(q34;q11.2); BCR-ABL1
CL374485|T191|Philadelphia Positive Childhood Precursor Lymphoblastic Leukemia
CL374485|T191|Philadelphia Positive Childhood Acute Lymphoblastic Leukemia
C1706717|T049|Adenosine to Guanosine Transition Abnormality
C1706717|T049|Adenosine to Guanosine Transition
C1706717|T049|Adenosine to Guanosine Mutation
C0742352|T033|Chest Wall Mass
C0742352|T033|Chest wall mass
C0742352|T033|Chest mass NOS
C0742352|T033|Chest Mass
C0742352|T033|Chest mass
C0742352|T033|CHEST MASS
C0742352|T033|chest mass
C0742352|T033|Mass of chest wall (finding)
C0742352|T033|thoracic mass
C0742352|T033|Mass of chest wall
C0684830|T191|Metastatic Malignant Neoplasm to the Axilla
C0684830|T191|Axillary Metastases
C0684830|T191|Metastatic Malignant Tumor to the Axilla
C0684830|T191|Axillary Metastasis
CL472832|T191|Recurrent Malignant Extragonadal Non-Seminomatous Germ Cell Tumor
C0221286|T191|Paget Disease of the Penis
C0221286|T191|Paget's Disease of Penis
C0221286|T191|Penile adenocarcinoma
C0221286|T191|Paget's Disease of the Penis
C1334037|T191|Classical Hodgkin Lymphoma Type Post-Transplant Lymphoproliferative Disorder
C1334037|T191|Hodgkin Lymphoma Post-Transplant Lymphoproliferative Disorder
C1334037|T191|Hodgkin's Lymphoma Post-Transplant Lymphoproliferative Disorder
C1334037|T191|Classical Hodgkin Lymphoma Type PTLD
C1334037|T191|Hodgkin Lymphoma PTLD
C1334037|T191|Classical Hodgkin Lymphoma Post-Transplant Lymphoproliferative Disorder
C1334037|T191|Hodgkin's Lymphoma PTLD
C0280367|T191|Recurrent Oral Cavity Adenoid Cystic Carcinoma
C0280367|T191|Relapsed Oral Cavity Adenoid Cystic Carcinoma
C0280367|T191|Recurrent Mouth Adenoid Cystic Carcinoma
C0280367|T191|adenoid cystic carcinoma of the oral cavity, recurrent
C0280367|T191|recurrent adenoid cystic carcinoma of the oral cavity
C0280367|T191|Relapsed Adenoid Cystic Carcinoma of Mouth
C0280367|T191|oral cavity adenoid cystic carcinoma, recurrent
C0280367|T191|Recurrent Adenoid Cystic Carcinoma of Oral Cavity
C0280367|T191|Relapsed Adenoid Cystic Carcinoma of the Oral Cavity
C0280367|T191|Relapsed Adenoid Cystic Carcinoma of Oral Cavity
C0280367|T191|Adenoid cystic carcinoma of the oral cavity recurrent
C0280367|T191|Recurrent Adenoid Cystic Carcinoma of the Oral Cavity
C0280367|T191|Relapsed Adenoid Cystic Carcinoma of the Mouth
C0280367|T191|Recurrent Adenoid Cystic Carcinoma of the Mouth
C0280367|T191|Recurrent Adenoid Cystic Carcinoma of Mouth
C0280367|T191|Relapsed Mouth Adenoid Cystic Carcinoma
C1304517|T191|Extrarenal Rhabdoid Tumor
C1304517|T191|Malignant Extrarenal Rhabdoid Neoplasm
C1304517|T191|Extrarenal rhabdoid tumor (disorder)
C1304517|T191|Extrarenal rhabdoid tumour
C1304517|T191|Extrarenal rhabdoid tumor
C0685943|T191|Metastatic Malignant Neoplasm to the Lip
C0685943|T191|Metastasis to the Lip
C0685943|T191|Metastatic Tumor to the Lip
C0685943|T191|Metastatic Neoplasm to the Lip
C0441959|T033|Node stage N0
C0441959|T033|N0 Stage
C0441959|T033|N0 category (finding)
C0441959|T033|N0 TNM Finding
C0441959|T033|N0 Regional Lymph Nodes Finding
C0441959|T033|N0 Lymph Node Stage
C0441959|T033|N0 category
C0441959|T033|N0 Cancer Stage Finding
C0441959|T033|N0 Node Finding
C0441959|T033|Lymph Node Stage N0
C0441959|T033|N0 Stage Finding
C0441959|T033|N0
C0441959|T033|Node Stage N0
C0441959|T033|N0 Lymph Node Finding
C0441959|T033|N0 lymph node stage
C0441959|T033|N0 stage
C0441959|T033|N0 Regional Lymph Node Stage Finding
C0441959|T033|N0 Node Stage
C0730492|T170|Tumor stage Tis pu
C0730492|T170|Tumor stage Tis pu (finding)
C0730492|T170|Tumour stage Tis pu
C1518870|T191|Pancreatic Mucinous-Cystic Neoplasm with an Associated Invasive Carcinoma
C1518870|T191|Pancreatic Invasive Mucinous Cystadenocarcinoma
C1518870|T191|Pancreatic Mucinous Cystic Neoplasm with an Associated Invasive Carcinoma
C2347915|T191|Recurrent Grade III Lymphomatoid Granulomatosis
C1517281|T061|Focused Ultrasound Therapy
C1517281|T061|Therapy (Focused US)
C1517281|T061|Therapy, Focused Ultrasound
C1517281|T061|Focused Ultrasound
C1517281|T061|High Power Focused Ultrasound
C1512363|T061|Helium-Ion Radiation
C0278700|T191|Recurrent Childhood Liver Cancer
C0278700|T191|Relapsed Pediatric Cancer of the Liver
C0278700|T191|Recurrent Childhood Cancer of Liver
C0278700|T191|pediatric liver cancer, recurrent
C0278700|T191|Recurrent Pediatric Cancer of Liver
C0278700|T191|Relapsed Pediatric Liver Cancer
C0278700|T191|Recurrent Pediatric Cancer of the Liver
C0278700|T191|recurrent childhood liver cancer
C0278700|T191|Recurrent Childhood Cancer of the Liver
C0278700|T191|Relapsed Childhood Liver Cancer
C0278700|T191|liver cancer, childhood, recurrent
C0278700|T191|Relapsed Childhood Cancer of Liver
C0278700|T191|Relapsed Childhood Cancer of the Liver
C0278700|T191|Recurrent Pediatric Liver Cancer
C0278700|T191|liver cancer, pediatric, recurrent
C0278700|T191|Relapsed Pediatric Cancer of Liver
C0278700|T191|childhood liver cancer, recurrent
C0278700|T191|recurrent pediatric liver cancer
C1384494|T191|Secondary Carcinoma
C1384494|T191|Carcinoma, metastatic, NOS
C1384494|T191|Metastatic carcinoma
C1384494|T191|Secondary carcinoma
C1384494|T191|Carcinoma, metastatic
C1384494|T191|Metastatic Carcinoma
C1384494|T191|Carcinoma, metastatic (morphologic abnormality)
C1384494|T191|METASTATIC CARCINOMA
C0220644|T191|Childhood Hodgkin Lymphoma
C0220644|T191|childhood Hodgkin disease
C0220644|T191|Childhood HD
C0220644|T191|Hodgkin's disease, childhood
C0220644|T191|Pediatric Hodgkin's Disease
C0220644|T191|Hodgkin lymphoma, child
C0220644|T191|Childhood Hodgkin's Lymphoma
C0220644|T191|Childhood Hodgkin's Disease
C0220644|T191|HD, childhood
C0220644|T191|childhood Hodgkin lymphoma
C0220644|T191|lymphoma, Hodgkin's, childhood
C0220644|T191|Pediatric Hodgkin's Lymphoma
C0220644|T191|pediatric HD
C0220644|T191|childhood Hodgkins disease
C0220644|T191|Pediatric HD
C0220644|T191|childhood HD
C0220644|T191|Lymphoma, Hodgkin lymphoma, child
C0220644|T191|childhood Hodgkin's disease
C0220644|T191|Hodgkin's lymphoma, childhood
C0220644|T191|pediatric Hodgkin's disease
C0220644|T191|childhood Hodgkin's lymphoma
C0220644|T191|childhood Hodgkins lymphoma
C0346974|T191|Metastatic Malignant Neoplasm to the Colon
C0346974|T191|Metastatic Neoplasm to the Colon
C0346974|T191|Metastatic Tumor to the Colon
C1524020|T061|Radiation Ionizing Radiotherapy
C1524020|T061|Radiation
C0278952|T191|Recurrent Nasopharynx Carcinoma
C0278952|T191|Recurrent Carcinoma of the Nasopharynx
C0278952|T191|Recurrent Cancer of Nasopharynx
C0278952|T191|Relapsed Cancer of Nasopharynx
C0278952|T191|Relapsed Nasopharynx Carcinoma
C0278952|T191|Relapsed Cancer of the Nasopharynx
C0278952|T191|Relapsed Nasopharyngeal Cancer
C0278952|T191|Relapsed Nasopharyngeal Carcinoma
C0278952|T191|nasopharynx cancer, recurrent
C0278952|T191|Nasopharyngeal cancer recurrent
C0278952|T191|Recurrent Carcinoma of Nasopharynx
C0278952|T191|Relapsed Carcinoma of the Nasopharynx
C0278952|T191|Recurrent Nasopharyngeal Cancer
C0278952|T191|Nasopharyngeal Cancer, Recurrent
C0278952|T191|recurrent nasopharyngeal cancer
C0278952|T191|Relapsed Carcinoma of Nasopharynx
C0278952|T191|Recurrent Cancer of the Nasopharynx
C0278952|T191|Recurrent Nasopharyngeal Carcinoma
C0278952|T191|nasopharyngeal cancer, recurrent
C1334807|T191|Mucinous Breast Carcinoma
C1334807|T191|Invasive Mucinous Breast Carcinoma
C1334807|T191|Mucinous Carcinoma of Breast
C1334807|T191|ductal mucinous breast carcinoma
C1334807|T191|Mucinous carcinoma of breast
C1334807|T191|Mucinous ductal breast carcinoma
C1334807|T191|Colloid Carcinoma of Breast
C1334807|T191|Colloid Breast Carcinoma
C1334807|T191|colloid ductal breast carcinoma
C1334807|T191|Infiltrating Mucinous Breast Carcinoma
C1334807|T191|Colloid Carcinoma of the Breast
C1334807|T191|Invasive Colloid Breast Carcinoma
C1334807|T191|Mucinous Carcinoma of the Breast
C1334807|T191|Mucinous carcinoma of breast (disorder)
C1334807|T191|Breast Mucinous Carcinoma
C1334807|T191|Infiltrating Colloid Breast Carcinoma
C1334807|T191|ductal colloid breast carcinoma
C1334807|T191|mucinous ductal breast carcinoma
C1334807|T191|Mucinous breast carcinoma
C0877357|T191|Recurrent Gallbladder Carcinoma
C0877357|T191|Recurrent Gallbladder Cancer
C0877357|T191|Gallbladder cancer recurrent
C0877357|T191|Recurrent Cancer of the Gallbladder
C0877357|T191|Recurrent Cancer of Gallbladder
C0877357|T191|Relapsed Cancer of the Gallbladder
C0877357|T191|Malignant neoplasm of gallbladder recurrent
C0877357|T191|Gallbladder carcinoma recurrent
C0877357|T191|recurrent gallbladder cancer
C0877357|T191|Relapsed Gallbladder Cancer
C0877357|T191|gallbladder cancer, recurrent
C0877357|T191|Gallbladder Cancer, Recurrent
C0877357|T191|Relapsed Cancer of Gallbladder
C1883258|T061|TCH Regimen
C1883258|T061|Docetaxel-Carboplatin-Trastuzumab Regimen
C1883258|T061|Taxotere-Carboplatin-Herceptin Regimen
C0240007|T033|Inguinal Mass
C0240007|T033|Inguinal mass
C0240007|T033|Groin mass
C0240007|T033|Groin mass (finding)
C0240007|T033|INGUINAL MASS
C0240007|T033|Groin lump
C0240007|T033|Mass of inguinal region
C0475384|T185|Tumor stage T1a2
C0475384|T185|Tumour stage T1a2
C0475384|T185|Tumor stage T1a2 (finding)
C0278699|T191|Stage IV Childhood Hepatocellular Carcinoma
C0278699|T191|Stage IV Pediatric Hepatoma
C0278699|T191|Stage IV Childhood Hepatocellular Carcinoma AJCC v7
C0278699|T191|Stage IV Pediatric Hepatocellular Carcinoma
C0278699|T191|Stage IV Pediatric Liver Cell Carcinoma
C0278699|T191|Stage IV Childhood Hepatoma
C0278699|T191|stage IV childhood liver cancer
C0278699|T191|Stage IV Childhood Liver Cell Carcinoma
C1332989|T191|Childhood Ovarian Embryonal Carcinoma
C1332989|T191|Childhood Embryonal Carcinoma of Ovary
C1332989|T191|Pediatric Embryonal Carcinoma of the Ovary
C1332989|T191|Pediatric Ovarian Embryonal Carcinoma
C1332989|T191|Pediatric Embryonal Carcinoma of Ovary
C1332989|T191|Childhood Embryonal Carcinoma of the Ovary
C1332948|T191|Childhood Brain Germinoma
C1332948|T191|Germinoma of the Pediatric Brain
C1332948|T191|Pediatric Brain Germ Cell Cancer
C1332948|T191|Pediatric Brain Germinoma
C1332948|T191|Germinoma of Pediatric Brain
C1332948|T191|Germinoma of the Childhood Brain
C1332948|T191|Germinoma of Childhood Brain
C1333313|T191|Drop Metastasis to Spinal Cord
C1333313|T191|Drop Metastatic Tumor to the Spinal Cord
C1333313|T191|Drop Secondary Malignant Tumor to the Spinal Cord
C1333313|T191|Drop Secondary Malignant Neoplasm to the Spinal Cord
C1333313|T191|Drop Metastatic Neoplasm to the Spinal Cord
C0563528|T061|Right Oophorectomy
C0563528|T061|Oophorectomy right
C0563528|T061|Right oophorectomy
C0563528|T061|Right oophorectomy (procedure)
C0279943|T191|Recurrent Childhood Soft Tissue Sarcoma
C0279943|T191|recurrent childhood soft tissue sarcoma
C0279943|T191|Recurrent Childhood Sarcoma of the Soft Tissue
C0279943|T191|STS, childhood, recurrent
C0279943|T191|Relapsed Pediatric Sarcoma of the Soft Tissue
C0279943|T191|pediatric soft tissue sarcoma, recurrent
C0279943|T191|Relapsed Pediatric Soft Tissue Sarcoma
C0279943|T191|Relapsed Childhood Sarcoma of the Soft Tissue
C0279943|T191|Recurrent Pediatric Soft Tissue Sarcoma
C0279943|T191|childhood STS, recurrent
C0279943|T191|Recurrent Pediatric Sarcoma of the Soft Tissue
C0279943|T191|Recurrent Childhood Sarcoma of Soft Tissue
C0279943|T191|pediatric STS, recurrent
C0279943|T191|Relapsed Childhood Sarcoma of Soft Tissue
C0279943|T191|childhood soft tissue sarcoma, recurrent
C0279943|T191|STS, recurrent, childhood
C0279943|T191|Relapsed Childhood Soft Tissue Sarcoma
C0279943|T191|Relapsed Pediatric Sarcoma of Soft Tissue
C0279943|T191|Recurrent Pediatric Sarcoma of Soft Tissue
C0475400|T185|Tumor stage T1a1
C0475400|T185|Tumor stage T1a1 (finding)
C0475400|T185|Tumour stage T1a1
C0279754|T034|Estrogen Receptor Positive
C0279754|T034|positive estrogen receptor
C0279754|T034|estrogen receptor positive
C0279754|T034|Positive Estrogen Receptor
C0279754|T034|ER+
C3272449|T033|N1bII Stage Finding
C0855045|T191|Recurrent Extraosseous Ewing Sarcoma
C0855045|T191|Recurrent Extra-Osseous Ewing's Sarcoma
C0855045|T191|Extra-osseous Ewing's sarcoma recurrent
C0855045|T191|Recurrent Extraosseous Ewing's Sarcoma
C0855045|T191|Extra-Osseous Ewing's Sarcoma, Recurrent
C0855045|T191|Relapsed Extra-Osseous Ewing's Sarcoma
C0855045|T191|Recurrent Extraskeletal Ewing's Sarcoma
C0337666|T055|Cigar Smoking
C0337666|T055|Cigar Smokings
C0337666|T055|Smoking, Cigar
C0337666|T055|Cigar smoker (finding)
C0337666|T055|Cigar smoking
C0337666|T055|Smokings, Cigar
C0337666|T055|Cigar smoker
C1335256|T191|PRETEXT Stage 2 Hepatoblastoma
C1333126|T033|Comedo-Like Necrosis
C0029189|T061|Orchiectomy
C0029189|T061|Total orchidectomy (procedure)
C0029189|T061|orchidectomy
C0029189|T061|Orchidectomies
C0029189|T061|Orchiectomies
C0029189|T061|Testis excision (procedure)
C0029189|T061|Orchidectomy
C0029189|T061|Orchidectomy NOS
C0029189|T061|ORCHIECTOMY
C0029189|T061|Excision of testis
C0029189|T061|male gonadectomy
C0029189|T061|Male Gonadectomy
C0029189|T061|Testis excision
C0029189|T061|Castration
C0029189|T061|Male Castration
C0029189|T061|Total orchidectomy
C0029189|T061|orchiectomy
C0346976|T191|Metastatic Malignant Neoplasm to the Pancreas
C0346976|T191|Secondary Malignant Neoplasm to the Pancreas
C0346976|T191|Secondary Malignant Tumor to the Pancreas
C0346976|T191|Metastatic Tumor to the Pancreas
C0346976|T191|Secondary Cancer to the Pancreas
C0346976|T191|Metastatic Cancer to the Pancreas
C0346976|T191|Metastatic Neoplasm to the Pancreas
C1335703|T191|Recurrent Head and Neck Carcinoma
C1335703|T191|Recurrent Head and Neck Cancer
C1332057|T191|AIDS-Related Plasmablastic Lymphoma of the Oral Mucosa
C1332057|T191|AIDS-Related Plasmablastic Lymphoma of Oral Mucosa
C0279916|T191|Stage III Childhood Hodgkin Lymphoma
C0279916|T191|Childhood Hodgkin's Disease Stage III
C0279916|T191|Pediatric Hodgkin's Lymphoma Stage III
C0279916|T191|Stage III Pediatric Hodgkin's Lymphoma
C0279916|T191|Childhood Hodgkin's Lymphoma Stage III
C0279916|T191|Stage III Childhood Hodgkin's Lymphoma
C0279916|T191|stage III childhood Hodgkin lymphoma
C0279916|T191|Pediatric Hodgkin's Disease Stage III
C0424864|T033|Width of lump
C0424864|T033|Width of lump (observable entity)
C0424864|T033|Breadth of lump
C1332962|T191|Childhood Cerebral Ependymoblastoma
C1332962|T191|Pediatric Cerebral Ependymoblastoma
C0730493|T170|Tumor stage Tis pd
C0730493|T170|Tumor stage Tis pd (finding)
C0730493|T170|Tumour stage Tis pd
C1334748|T191|Methotrexate-Associated Hodgkin Lymphoma
C1334748|T191|Methotrexate-Associated Hodgkin's Lymphoma
C1511302|T191|Breast Carcinoma with Choriocarcinomatous Features
C0153678|T191|Metastatic Malignant Neoplasm to the Pleura
C0153678|T191|Metastatic Tumor to the Pleura
C0153678|T191|Metastatic Neoplasm to the Pleura
C0153678|T191|Metastases to Pleura
C0153678|T191|Metastasis to the Pleura
C1377604|T191|Childhood Central Nervous System Choriocarcinoma
C1377604|T191|Choriocarcinoma of Pediatric Central Nervous System
C1377604|T191|Choriocarcinoma of the Pediatric CNS
C1377604|T191|Choriocarcinoma of the Pediatric Central Nervous System
C1377604|T191|Choriocarcinoma of Childhood Central Nervous System
C1377604|T191|childhood CNS choriocarcinoma
C1377604|T191|Childhood CNS Choriocarcinoma
C1377604|T191|Pediatric Central Nervous System Choriocarcinoma
C1377604|T191|Choriocarcinoma of the Childhood CNS
C1377604|T191|Choriocarcinoma of the Childhood Central Nervous System
C1377604|T191|Pediatric CNS Choriocarcinoma
C1377604|T191|Choriocarcinoma of Pediatric CNS
C1377604|T191|Choriocarcinoma of Childhood CNS
C1377604|T191|childhood central nervous system choriocarcinoma
C1332048|T191|AIDS-Related Large B-Cell Lymphoma Arising in Human Herpes Virus 8-Associated Multicentric Castleman Disease
C1332048|T191|AIDS-Related Kaposi Sarcoma-Associated Human Herpes Virus 8 Positive Extracavity Lymphoma
C1332048|T191|AIDS-Related Kaposi's Sarcoma-Associated Human Herpes Virus 8 Positive Extracavity Lymphoma
C1332048|T191|AIDS-Related Large B-Cell Lymphoma Arising in HHV 8-Associated Multicentric Castleman Disease
C1335446|T191|Poorly Differentiated Prostate Adenocarcinoma
C2825187|T061|Septal Ablation
C2825187|T061|SEPTAL ABLATION
C1334044|T033|Hormone Responsive Mass
C1321208|T033|Tumor size, right ovary
C1321208|T033|Tumor size, right ovary (observable entity)
C1321208|T033|Tumour size, right ovary
C1332039|T191|AIDS-Related Carcinoma
C1332039|T191|AIDS Related Carcinoma
C0854755|T191|Recurrent Lip and Oral Cavity Carcinoma
C0854755|T191|Recurrent Lip and Oral Cavity Cancer
C2986603|T061|Intraperitoneal Radiation Therapy
C2986603|T061|intraperitoneal radiation therapy
C1512710|T045|Induced Mutation
C1512710|T045|induced_mutation
C1512710|T045|Induced DNA Alteration
C1512710|T045|Induced Sequence Alteration
C0475389|T185|T2c Stage Finding
C0475389|T185|T2c TNM Finding
C0475389|T185|T2c Stage
C0475389|T185|T2c Tumor Finding
C0475389|T185|T2c Tumor Stage
C0475389|T185|Tumor stage T2c (finding)
C0475389|T185|T2c Primary Tumor Finding
C0475389|T185|Tumor stage T2c
C0475389|T185|T2c
C0475389|T185|Tumour stage T2c
C0475389|T185|T2c Cancer Stage Finding
C0475389|T185|Tumor Stage T2c
C0475389|T185|T2c Primary Tumor Stage Finding
C0730459|T170|Tumor stage T1b2
C0730459|T170|Tumor stage T1b2 (finding)
C0730459|T170|Tumour stage T1b2
C0279613|T191|Childhood Alveolar Rhabdomyosarcoma
C0279613|T191|Alveolar Childhood Rhabdomyosarcoma
C0279613|T191|alveolar childhood rhabdomyosarcoma
C0279613|T191|Pediatric Alveolar Rhabdomyosarcoma
C0279613|T191|alveolar pediatric rhabdomyosarcoma
C0279613|T191|childhood rhabdomyosarcoma, alveolar
C0279613|T191|rhabdomyosarcoma, pediatric alveolar
C0279613|T191|pediatric rhabdomyosarcoma, alveolar
C0279613|T191|rhabdomyosarcoma, alveolar childhood
C0279613|T191|rhabdomyosarcoma, childhood alveolar
C0730458|T170|Tumor stage T1b1
C0730458|T170|Tumor stage T1b1 (finding)
C0730458|T170|Tumour stage T1b1
C1337020|T191|Well Differentiated Prostate Adenocarcinoma
CL033795|T191|Recurrent Nasal Cavity and Paranasal Sinus Carcinoma
CL033795|T191|Recurrent Nasal Cavity and Paranasal Sinus Cancer
C2347757|T191|Childhood Classical Hodgkin Lymphoma
C116431|T061|Active Breathing Coordinator-Mediated Radiation Therapy
C116431|T061|ABC
C116431|T061|Active Breathing Coordinator
C1332956|T191|Childhood Central Nervous System Mixed Germ Cell Tumor
C1332956|T191|childhood central nervous system mixed germ cell tumor
C1332956|T191|childhood CNS mixed germ cell tumor
C1336022|T191|Solar Radiation-Related Malignant Neoplasm
C1336022|T191|Solar Radiation-Related Cancer
C1336835|T049|Tumor Cell Necrosis
CL448519|T191|Recurrent Salivary Gland Carcinoma
CL448519|T191|recurrent salivary gland cancer
CL448519|T191|Recurrent Cancer of Salivary Gland
CL448519|T191|Relapsed Carcinoma of Salivary Gland
CL448519|T191|Relapsed Cancer of Salivary Gland
CL448519|T191|Recurrent Cancer of the Salivary Gland
CL448519|T191|Recurrent Carcinoma of the Salivary Gland
CL448519|T191|Recurrent Carcinoma of Salivary Gland
CL448519|T191|Relapsed Cancer of the Salivary Gland
CL448519|T191|Relapsed Salivary Gland Cancer
CL448519|T191|Relapsed Carcinoma of the Salivary Gland
CL448519|T191|Recurrent Salivary Gland Cancer
CL448519|T191|Salivary Gland Cancer, Recurrent
CL448519|T191|salivary gland cancer, recurrent
CL448519|T191|Relapsed Salivary Gland Carcinoma
C0441917|T033|L0 Stage Finding
C0441917|T033|L0 TNM Finding
C0441917|T033|Lymphatic stage L0
C0441917|T033|L0 Stage
C0441917|T033|L0 Cancer Stage Finding
C0441917|T033|Lymphatic Stage L0
C0441917|T033|L0
C0441917|T033|L0 stage (finding)
C0441917|T033|L0 Lymphatic Vessel Invasion Finding
C0441917|T033|L0 Lymphatic Invasion Finding
C0441917|T033|L0 stage
C0441917|T033|L0 Lymphatic Stage
C0441917|T033|L0: no lymphatic vessel invasion
C1335503|T191|Prostate Adenosquamous Carcinoma
C1335503|T191|Adenosquamous Carcinoma of the Prostate
C1335503|T191|Adenosquamous Carcinoma of Prostate
C1334717|T191|Metastatic Carcinoma to the Adrenal Medulla
C1334717|T191|Metastatic Carcinoma to Adrenal Medulla
C1334717|T191|Adrenal Medulla Carcinoma
C1332038|T191|AIDS-Related Anal Carcinoma
C1332038|T191|AIDS-related anal cancer
C1332038|T191|AIDS-Related Anal Cancer
C0334373|T191|Infiltrating Papillary Adenocarcinoma
C0334373|T191|Infiltrating and papillary adenocarcinoma
C0334373|T191|Intraductal papillary adenocarcinoma with invasion
C0334373|T191|Intraductal papillary adenocarcinoma with invasion (morphologic abnormality)
C0334373|T191|[M]Intraductal papillary adenocarcinoma with invasion
C0334373|T191|Infiltrating papillary adenocarcinoma
C0334373|T191|Intraductal Papillary Adenocarcinoma with Invasion
C0334373|T191|[M] Intraductal papillary adenocarcinoma with invasion
C1880765|T033|Fetiform Mass
C1880881|T061|GT Regimen
C1880881|T061|Gemcitabine-Taxol Regimen
C0280787|T191|Adult Anaplastic Ependymoma
C0280787|T191|anaplastic ependymoma, adult
C0280787|T191|adult malignant ependymoma
C0280787|T191|Adult Malignant Ependymoma
C0280787|T191|malignant ependymoma, adult
C0280787|T191|adult anaplastic ependymoma
C0280787|T191|ependymoma, adult malignant
C0280787|T191|Malignant Adult Ependymoma
C0441962|T033|N1 Stage Finding
C0441962|T033|Node Stage N1
C0441962|T033|N1 TNM Finding
C0441962|T033|N1 category
C0441962|T033|N1 lymph node stage
C0441962|T033|N1 Stage
C0441962|T033|N1 Regional Lymph Nodes Finding
C0441962|T033|N1 category (finding)
C0441962|T033|N1 Lymph Node Finding
C0441962|T033|Node stage N1
C0441962|T033|N1 Cancer Stage Finding
C0441962|T033|N1 Regional Lymph Node Stage Finding
C0441962|T033|N1 stage
C0441962|T033|N1 Node Finding
C0441962|T033|N1 Node Stage
C0441962|T033|N1
C0441962|T033|N1 Lymph Node Stage
C0441962|T033|Lymph Node Stage N1
C1519559|T061|Total Estrogen Blockade
C1519559|T061|total estrogen blockade
C0441918|T033|L1 stage
C0441918|T033|L1 Lymphatic Invasion Finding
C0441918|T033|L1: lymphatic vessel invasion
C0441918|T033|L1 Stage
C0441918|T033|L1 Lymphatic Stage
C0441918|T033|L1 TNM Finding
C0441918|T033|L1 Lymphatic Vessel Invasion Finding
C0441918|T033|L1 Stage Finding
C0441918|T033|L1 Cancer Stage Finding
C0441918|T033|Lymphatic stage L1
C0441918|T033|Lymphatic Stage L1
C0441918|T033|L1 stage (finding)
C0441918|T033|L1
C0220645|T191|Childhood Soft Tissue Sarcoma
C0220645|T191|Pediatric Sarcoma of Soft Tissue
C0220645|T191|Pediatric Sarcoma of the Soft Tissue
C0220645|T191|Childhood Sarcoma of the Soft Tissue
C0220645|T191|childhood soft tissue sarcoma
C0220645|T191|STS, childhood
C0220645|T191|soft tissue sarcoma, childhood
C0220645|T191|Childhood Sarcoma of Soft Tissue
C0220645|T191|Pediatric Soft Tissue Sarcoma
C0220645|T191|Soft tissue sarcoma, child
C0220645|T191|pediatric soft tissue sarcoma
C0220645|T191|pediatric STS
C0220645|T191|childhood STS
C0278878|T191|Adult Glioblastoma
C0278878|T191|grade IV adult astrocytoma
C0278878|T191|CNS tumor, adult grade IV astrocytoma
C0278878|T191|CNS tumor, grade IV adult astrocytoma
C0278878|T191|glioblastoma multiforme, adult
C0278878|T191|adult CNS tumor, glioblastoma multiforme
C0278878|T191|adult glioblastoma
C0278878|T191|Grade IV Adult Astrocytic Tumor
C0278878|T191|adult glioblastoma multiforme
C0278878|T191|astrocytoma, grade IV adult
C0278878|T191|glioblastoma, adult
C0278878|T191|Grade IV Adult Astrocytic Neoplasm
C0278878|T191|CNS tumor, adult glioblastoma multiforme
C0278878|T191|Adult Glioblastoma Multiforme
C0278878|T191|central nervous system tumor, astrocytoma, grade IV adult
C1333005|T191|Childhood Systemic Anaplastic Large Cell Lymphoma
C1333005|T191|Pediatric Systemic CD30+ Anaplastic Large Cell Lymphoma
C1333005|T191|Pediatric Systemic Anaplastic Large Cell Lymphoma
C1333005|T191|Childhood Systemic CD30+ Anaplastic Large Cell Lymphoma
C1333005|T191|Childhood Systemic K-1+ Anaplastic Large Cell Lymphoma
C1333005|T191|Pediatric Systemic K-1+ Anaplastic Large Cell Lymphoma
C1332128|T191|Peritoneal Carcinomatosis
C1332128|T191|Carcinomatosis of the Peritoneum
C1332128|T191|Peritoneal carcinomatosis
C1332128|T191|Abdominal Carcinomatosis
C1332128|T191|peritoneal carcinomatosis
C0153676|T191|Metastatic Malignant Neoplasm to the Lung
C0153676|T191|Metastatic Tumor to the Lung
C0153676|T191|Metastasis to Lung
C0153676|T191|Metastases to lung, NOS
C0153676|T191|Metastases to Lung
C0153676|T191|Metastasis to the Lung
C0153676|T191|Lung Metastases
C0153676|T191|Metastatic Neoplasm to the Lung
C0153676|T191|lung metastasis
C1707606|T049|Cytosine to Thymidine Transition Abnormality
C1707606|T049|Cytosine to Thymidine Mutation
C1707606|T049|Cytosine to Thymidine Transition
C0886477|T191|Childhood Malignant Testicular Germ Cell Tumor
C0886477|T191|Childhood Testicular Germ Cell Neoplasm
C0886477|T191|pediatric testicular germ cell tumor
C0886477|T191|childhood testicular germ cell tumor
C0886477|T191|Pediatric Testicular Germ Cell Tumor
C0886477|T191|testicular germ cell tumor, pediatric
C0886477|T191|germ cell tumor, testicular, childhood
C0886477|T191|germ cell tumor, testicular, pediatric
C0886477|T191|Pediatric Testicular Germ Cell Neoplasm
C0886477|T191|testicular germ cell tumor, childhood
C0886477|T191|childhood malignant testicular germ cell tumor
C0886477|T191|Childhood Testicular Germ Cell Tumor
C0240611|T033|Ovarian Mass
C0240611|T033|Ovarian mass
C0240611|T033|Mass of ovary
C0240611|T033|OVARIAN MASS
C0240611|T033|Mass of Ovary
C0240611|T033|Mass of ovary (finding)
C1833921|T191|Hereditary Thyroid Gland Medullary Carcinoma
C1833921|T191|Familial medullary thyroid carcinoma
C1833921|T191|THYROID CARCINOMA, FAMILIAL MEDULLARY
C1833921|T191|familial medullary thyroid cancer
C1833921|T191|MTC
C1833921|T191|hereditary medullary thyroid cancer
C1833921|T191|Medullary thyroid cancer, familial
C1833921|T191|MTC1
C1833921|T191|Familial Thyroid Gland Medullary Carcinoma
C1833921|T191|hereditary thyroid gland medullary carcinoma
C1833921|T191|FMTC
C1833921|T191|Thyroid Carcinoma, Familial Medullary
C1833921|T191|familial thyroid gland medullary carcinoma
C1833921|T191|Thyroid cancer, familial medullary
C1833921|T191|Familial medullary thyroid cancer
CL034604|T191|Childhood Extragonadal Malignant Germ Cell Tumor
CL034604|T191|childhood extragonadal germ cell tumor
CL034604|T191|pediatric extragonadal germ cell tumor
CL034604|T191|germ cell tumor, extragonadal, childhood
CL034604|T191|extragonadal germ cell tumor, childhood
CL034604|T191|germ cell tumor, extragonadal, pediatric
CL034604|T191|extragonadal germ cell tumor, pediatric
C0206076|T201|Reproductive History
C0206076|T201|Histories, Reproductive
C0206076|T201|Reproductive Issues
C0206076|T201|History, Reproductive
C0206076|T201|reproductive issues
C0206076|T201|REPRODUCTIVE HIST
C0206076|T201|HIST REPRODUCTIVE
C0206076|T201|Reproductive Histories
C0206076|T201|Reproductive Factors
C0238729|T033|Axillary Mass
C0238729|T033|Axillary lump
C0238729|T033|Mass of axilla (finding)
C0238729|T033|Axillary mass
C0238729|T033|Lump of axilla
C0238729|T033|Mass of axilla
C0238729|T033|AXILLARY MASS
CL447332|T061|Fletcher-suit Brachytherapy
C0419095|T061|External Beam Radiation Therapy
C0419095|T061|Definitive Radiation Therapy
C0419095|T061|external radiation
C0419095|T061|Teletherapy
C0419095|T061|External beam radiotherapy
C0419095|T061|External Beam RT
C0419095|T061|external-beam radiation
C0419095|T061|Teleradiotherapy procedure (procedure)
C0419095|T061|External Radiation Therapy
C0419095|T061|EBRT
C0419095|T061|EB - External beam radiotherapy
C0419095|T061|Teletherapy procedure
C0419095|T061|external beam radiation therapy
C0419095|T061|Teleradiotherapy procedure
C0419095|T061|External Beam Radiotherapy
C0279922|T191|Childhood Mixed Cellularity Classical Hodgkin Lymphoma
C0279922|T191|Childhood Mixed Cellularity Hodgkin Lymphoma
C0279922|T191|mixed cellularity HD, childhood
C0279922|T191|pediatric Hodgkin's disease, mixed cellularity
C0279922|T191|Childhood Mixed Cellularity Hodgkin's Disease
C0279922|T191|lymphoma, mixed cellularity childhood Hodgkin's
C0279922|T191|mixed cellularity Hodgkin's disease, childhood
C0279922|T191|childhood mixed cellularity Hodgkin lymphoma
C0279922|T191|HD, mixed cellularity, childhood
C0279922|T191|MC HD, childhood
C0279922|T191|Hodgkin's disease, mixed cellularity, childhood
C0279922|T191|Pediatric MCHD
C0279922|T191|mixed cellularity childhood Hodgkin's disease
C0279922|T191|Childhood Mixed Cellularity Hodgkin's Lymphoma
C0279922|T191|childhood mixed cellularity Hodgkin's disease
C0279922|T191|MCHD, childhood
C0279922|T191|Pediatric Mixed Cellularity Hodgkin's Disease
C0279922|T191|pediatric mixed cellularity Hodgkin's disease
C0279922|T191|childhood Hodgkin's disease, mixed cellularity
C0279922|T191|childhood HD, mixed cellularity
C0279922|T191|Childhood MCHD
C0279922|T191|pediatric HD, mixed cellularity
C0279922|T191|Pediatric Mixed Cellularity Hodgkin's Lymphoma
CL376152|T191|Childhood Unfavorable Prognosis Hodgkin Lymphoma
CL376152|T191|childhood unfavorable prognosis Hodgkin lymphoma
C0745390|T047|Intrauterine Mass
C0745390|T047|Mass of Uterine Corpus
C0745390|T047|Mass of Uterine Body
C0745390|T047|Uterine Body Mass
C0745390|T047|Uterine Corpus Mass
C0745390|T047|Mass of the Uterine Body
C0745390|T047|Mass of the Uterine Corpus
C1332979|T191|Childhood Lymphoma
C1332979|T191|Pediatric Lymphoma
C1879280|T191|Childhood Nasal Type Extranodal NK/T-Cell Lymphoma
C1332985|T191|Childhood Nodular Lymphocyte Predominant Hodgkin Lymphoma
C1332985|T191|childhood Hodgkin's disease, lymphocyte predominant
C1332985|T191|HD lymphocyte predominant, childhood
C1332985|T191|Childhood Nodular Lymphocyte Predominant Hodgkin's Lymphoma
C1332985|T191|pediatric HD, lymphocyte predominant
C1332985|T191|Pediatric Nodular Lymphocyte Predominant Hodgkin's Lymphoma
C1332985|T191|lymphocyte predominant Hodgkin's disease, childhood
C1332985|T191|childhood HD, lymphocyte predominant
C1332985|T191|Pediatric Nodular Lymphocyte Predominant Hodgkin's Disease
C1332985|T191|HDLP, childhood
C1332985|T191|lymphocyte predominant HD, childhood
C1332985|T191|Childhood Nodular Lymphocyte Predominant Hodgkin's Disease
C1332985|T191|lymphoma, lymphocyte predominant childhood Hodgkin's
C1332985|T191|Pediatric NLPHD
C1332985|T191|childhood lymphocyte predominant Hodgkin's disease
C1332985|T191|pediatric lymphocyte predominant Hodgkin's disease
C1332985|T191|Hodgkin's disease, lymphocyte predominant, childhood
C1332985|T191|childhood lymphocyte predominant Hodgkin lymphoma
C1332985|T191|LP HD, childhood
C1332985|T191|pediatric Hodgkin's disease, lymphocyte predominant
C1332985|T191|LPHD, childhood
C1332985|T191|Childhood NLPHD
C1332985|T191|HD LP, childhood
C1332985|T191|childhood nodular lymphocyte predominant Hodgkin lymphoma
C1335433|T191|Pleural Carcinomatosis
C1335433|T191|Carcinomatosis of the Pleura
C114831|T191|Metastatic Malignant Neoplasm to Soft Tissues
C1334556|T191|ACTH-Producing Pituitary Gland Carcinoma
C1334556|T191|Malignant Adrenocorticotropin Producing Neoplasm of Pituitary Gland
C1334556|T191|Malignant ACTH Secreting Tumor of Pituitary
C1334556|T191|Malignant Adrenocorticotropin Producing Neoplasm of Pituitary
C1334556|T191|Malignant ACTH Secreting Pituitary Tumor
C1334556|T191|Malignant Adrenocorticotropin Producing Neoplasm of the Pituitary Gland
C1334556|T191|Malignant Adrenocorticotropin Producing Tumor of Pituitary
C1334556|T191|Malignant ACTH Secreting Tumor of Pituitary Gland
C1334556|T191|Malignant Adrenocorticotropin Secreting Pituitary Tumor
C1334556|T191|Malignant Corticotropin Secreting Pituitary Gland Neoplasm
C1334556|T191|Malignant Adrenocorticotropin Secreting Pituitary Gland Tumor
C1334556|T191|Malignant ACTH Secreting Neoplasm of the Pituitary
C1334556|T191|Malignant ACTH Producing Neoplasm of Pituitary
C1334556|T191|Malignant Adrenocorticotropin Producing Pituitary Gland Neoplasm
C1334556|T191|Malignant Corticotropinoma of Pituitary
C1334556|T191|Malignant Adrenocorticotropin Producing Pituitary Gland Tumor
C1334556|T191|Malignant Adrenocorticotropin Producing Tumor of the Pituitary
C1334556|T191|Malignant ACTH Producing Tumor of Pituitary Gland
C1334556|T191|Malignant Pituitary Gland Corticotropinoma
C1334556|T191|Malignant ACTH Producing Tumor of Pituitary
C1334556|T191|Malignant ACTH Producing Tumor of the Pituitary
C1334556|T191|Malignant ACTH Secreting Neoplasm of the Pituitary Gland
C1334556|T191|Malignant ACTH Producing Tumor of the Pituitary Gland
C1334556|T191|Malignant Adrenocorticotropin Producing Pituitary Tumor
C1334556|T191|Malignant Adrenocorticotropin Secreting Pituitary Gland Neoplasm
C1334556|T191|Malignant ACTH Secreting Pituitary Gland Tumor
C1334556|T191|Malignant ACTH Producing Pituitary Gland Neoplasm
C1334556|T191|Malignant Adrenocorticotropin Producing Tumor of the Pituitary Gland
C1334556|T191|Malignant ACTH Producing Pituitary Neoplasm
C1334556|T191|ACTH Producing Pituitary Gland Carcinoma
C1334556|T191|Malignant ACTH Producing Neoplasm of the Pituitary Gland
C1334556|T191|Malignant ACTH Secreting Tumor of the Pituitary Gland
C1334556|T191|Malignant Adrenocorticotropin Producing Pituitary Neoplasm
C1334556|T191|Malignant Pituitary Corticotropinoma
C1334556|T191|Malignant Corticotropinoma of the Pituitary Gland
C1334556|T191|Malignant ACTH Secreting Neoplasm of Pituitary
C1334556|T191|Malignant ACTH Secreting Pituitary Neoplasm
C1334556|T191|Malignant ACTH Producing Neoplasm of Pituitary Gland
C1334556|T191|Malignant Adrenocorticotropin Producing Neoplasm of the Pituitary
C1334556|T191|Malignant Adrenocorticotropin Producing Tumor of Pituitary Gland
C1334556|T191|Malignant ACTH Secreting Neoplasm of Pituitary Gland
C1334556|T191|Malignant ACTH Producing Pituitary Tumor
C1334556|T191|Malignant Adrenocorticotropin Secreting Pituitary Neoplasm
C1334556|T191|Malignant Corticotropinoma of the Pituitary
C1334556|T191|Malignant ACTH Producing Neoplasm of the Pituitary
C1334556|T191|Malignant ACTH Secreting Tumor of the Pituitary
C1334556|T191|Malignant ACTH Producing Pituitary Gland Tumor
C1334556|T191|Malignant Corticotropinoma of Pituitary Gland
C1707042|T191|Breast Carcinoma with Chondroid Metaplasia
C1707042|T191|Breast Carcinoma with Cartilaginous Metaplasia
C1514711|T061|Low-LET Radiotherapy
C1514711|T061|Radiotherapy, Low Linear Energy Transfer
C1514711|T061|Radiotherapy, Low LET
CL448348|T191|Childhood Supratentorial Ependymoblastoma
CL448348|T191|supratentorial ependymoblastoma, childhood
CL448348|T191|childhood supratentorial ependymoblastoma
CL448348|T191|ependymoblastoma, childhood supratentorial
CL448348|T191|Pediatric Supratentorial Ependymoblastoma
C0010408|T061|Cryosurgery
C0010408|T061|Cryoablation - action (qualifier value)
C0010408|T061|Cryosurgery - action (qualifier value)
C0010408|T061|Cryosurgery (procedure)
C0010408|T061|Cryoablations
C0010408|T061|CRYOSURG
C0010408|T061|cryoablation
C0010408|T061|CRYOABLATION
C0010408|T061|Cryosurgeries
C0010408|T061|Cryosurgery - action
C0010408|T061|cryosurgical ablation
C0010408|T061|Cryocautery - action (qualifier value)
C0010408|T061|Cryocautery
C0010408|T061|cryosurgery
C0010408|T061|Cryoablation - action
C0010408|T061|Cryocautery - action
C0010408|T061|Cryodestruction
C0010408|T061|Cryoablation
C2985381|T061|Systemic Radiation Therapy
C2985381|T061|systemic radiation therapy
C1335716|T191|Recurrent Nodular Lymphocyte Predominant Hodgkin Lymphoma
C1335716|T191|Relapsed Nodular Lymphocyte Predominant Hodgkin's Lymphoma
C1335716|T191|Recurrent Nodular Lymphocyte Predominant Hodgkin's Lymphoma
C1335716|T191|Recurrent Nodular Lymphocyte Predominant Hodgkin's Disease
C1335716|T191|Relapsed Nodular Lymphocyte Predominant Hodgkin's Disease
C1333009|T191|Childhood Testicular Mixed Germ Cell Neoplasm
C1333009|T191|Pediatric Testicular Mixed Germ Cell Tumor
C1333009|T191|Childhood Testicular Mixed Germ Cell Tumor
C1333009|T191|Pediatric Testicular Mixed Germ Cell Neoplasm
C114775|T191|Childhood Cerebral Neuroblastoma
C114775|T191|neuroblastoma, cerebral, pediatric
C114775|T191|childhood cerebral neuroblastoma
C114775|T191|neuroblastoma, cerebral, childhood
C114775|T191|neuroblastoma, childhood cerebral
C114775|T191|cerebral neuroblastoma, childhood
C114775|T191|pediatric cerebral neuroblastoma
C114775|T191|cerebral neuroblastoma, pediatric
C114775|T191|neuroblastoma, pediatric cerebral
CL448460|T191|Recurrent Malignant Gastric Neoplasm
C1334614|T191|Prolactin-Producing Pituitary Gland Carcinoma
C1334614|T191|Malignant Prolactin Secreting Neoplasm of the Pituitary Gland
C1334614|T191|Malignant Prolactin Producing Tumor of Pituitary
C1334614|T191|Malignant Prolactin Producing Neoplasm of the Pituitary
C1334614|T191|Malignant Prolactin Producing Tumor
C1334614|T191|PRL Producing Pituitary Gland Carcinoma
C1334614|T191|Malignant Prolactin Producing Neoplasm of the Pituitary Gland
C1334614|T191|Malignant Prolactin Producing Pituitary Tumor
C1334614|T191|Malignant Prolactin Producing Pituitary Gland Neoplasm
C1334614|T191|Malignant Pituitary Prolactinoma
C1334614|T191|Malignant Prolactin Producing Tumor of the Pituitary
C1334614|T191|Malignant Prolactin Producing Pituitary Neoplasm
C1334614|T191|Malignant Pituitary Gland Prolactinoma
C1334614|T191|Malignant Prolactin Producing Neoplasm of Pituitary
C1334614|T191|Malignant Prolactin Secreting Tumor of Pituitary Gland
C1334614|T191|Malignant Prolactin Secreting Tumor of the Pituitary Gland
C1334614|T191|Malignant Prolactin Secreting Tumor of Pituitary
C1334614|T191|Malignant Prolactinoma
C1334614|T191|Malignant Prolactin Producing Tumor of Pituitary Gland
C1334614|T191|Malignant Prolactin Secreting Pituitary Gland Neoplasm
C1334614|T191|Malignant Prolactinoma of Pituitary Gland
C1334614|T191|Malignant Prolactin Secreting Neoplasm of the Pituitary
C1334614|T191|Malignant Prolactin Secreting Neoplasm of Pituitary
C1334614|T191|Malignant Prolactin Producing Tumor of the Pituitary Gland
C1334614|T191|Malignant Prolactin Secreting Neoplasm of Pituitary Gland
C1334614|T191|Prolactin Producing Pituitary Gland Carcinoma
C1334614|T191|Malignant Prolactin Producing Pituitary Gland Tumor
C1334614|T191|Malignant Prolactin Secreting Tumor of the Pituitary
C1334614|T191|Malignant Prolactin Secreting Pituitary Tumor
C1334614|T191|Malignant Prolactinoma of the Pituitary Gland
C1334614|T191|Malignant Prolactinoma of Pituitary
C1334614|T191|Malignant Prolactin Secreting Pituitary Gland Tumor
C1334614|T191|Malignant Prolactin Secreting Pituitary Neoplasm
C1334614|T191|Malignant Prolactin Producing Neoplasm of Pituitary Gland
C1334614|T191|Malignant Prolactinoma of the Pituitary
C1301091|T201|Height of tumor at cut edge, after sectioning
C1301091|T201|Height of tumor at cut edge, after sectioning (observable entity)
C1301091|T201|Height of tumour at cut edge, after sectioning
C2985560|T061|Transarterial Radioembolization
C2985560|T061|intra-arterial brachytherapy
C2985560|T061|Radioembolisation
C2985560|T061|Radioembolization
C2985560|T061|radioembolization
C2985560|T061|transarterial radioembolization
C0278493|T191|Recurrent Breast Carcinoma
C0278493|T191|Breast Cancer, Recurrent
C0278493|T191|Carcinoma breast recurrent
C0278493|T191|Breast carcinoma recurrent
C0278493|T191|Breast carcinoma NOS recurrent
C0278493|T191|recurrent breast cancer
C0278493|T191|breast cancer, recurrent
C0278493|T191|Recurrent Breast Cancer
C0278493|T191|Breast cancer NOS recurrent
C0278493|T191|Breast cancer recurrent
C1377613|T191|Childhood Central Nervous System Yolk Sac Tumor
C1377613|T191|childhood CNS yolk sac tumor
C1377613|T191|Pediatric Central Nervous System Yolk Sac Tumor
C1377613|T191|childhood central nervous system yolk sac tumor
C1377613|T191|Pediatric Central Nervous System Yolk Sac Neoplasm
C1377613|T191|Pediatric Central Nervous System Endodermal Sinus Tumor
C1377613|T191|Pediatric Central Nervous System Endodermal Sinus Neoplasm
C1377613|T191|Childhood Central Nervous System Endodermal Sinus Neoplasm
C1377613|T191|Childhood Central Nervous System Endodermal Sinus Tumor
C1377613|T191|childhood CNS endodermal sinus tumor
C1377613|T191|Childhood Central Nervous System Yolk Sac Neoplasm
C1512418|T191|Hereditary Fallopian Tube Carcinoma
C1512418|T191|Familial Fallopian Tube Carcinoma
C0280364|T191|Recurrent Lip Basal Cell Carcinoma
C0280364|T191|Relapsed Lip Basal Cell Carcinoma
C0280364|T191|Recurrent Basal Cell Carcinoma of the Lip
C0280364|T191|Relapsed Basal Cell Carcinoma of the Lip
C0280364|T191|Recurrent Basal Cell Carcinoma of Lip
C0280364|T191|recurrent basal cell carcinoma of the lip
C0280364|T191|Relapsed Basal Cell Carcinoma of Lip
C0280364|T191|basal cell carcinoma of the lip, recurrent
C0280364|T191|lip basal cell carcinoma, recurrent
C1332242|T191|Ameloblastic Carcinoma Derived From Odontogenic Cyst
C1332242|T191|Ameloblastic Carcinoma Ex Odontogenic Cyst
C1336880|T191|Infiltrating Ureter Urothelial Carcinoma with Glandular Differentiation
C1336880|T191|Transitional Cell Carcinoma of the Ureter with Glandular Differentiation
C1336880|T191|Ureteral Transitional Cell Carcinoma with Glandular Differentiation
C1336880|T191|Transitional Cell Carcinoma of Ureter with Glandular Differentiation
C0349672|T191|Prostate Ductal Adenocarcinoma
C0349672|T191|Endometrioid carcinoma of prostate (disorder)
C0349672|T191|Ductal Adenocarcinoma of the Prostate
C0349672|T191|Prostate Endometrioid Adenocarcinoma
C0349672|T191|Endometrioid Carcinoma of the Prostate
C0349672|T191|Endometrioid Adenocarcinoma of the Prostate
C0349672|T191|Prostatic Endometrioid Carcinoma
C0349672|T191|Prostate Endometrioid Carcinoma
C0349672|T191|Ductal Adenocarcinoma of Prostate
C0349672|T191|Endometrioid carcinoma of prostate
C0349672|T191|Endometrioid Adenocarcinoma of Prostate
C0349672|T191|Endometrioid Carcinoma of Prostate
C0153690|T191|Metastatic Malignant Neoplasm to the Bone
C0153690|T191|Bone Metastases
C0153690|T191|Bone Metastasis
C0153690|T191|Metastatic Tumor to the Bone
C0153690|T191|Metastases to bone, NOS
C0153690|T191|Metastatic Cancer to the Bone
C0153690|T191|bone metastasis
C0153690|T191|Metastatic Neoplasm to the Bone
C1515865|T191|Acinar Prostate Adenocarcinoma, Oncocytic Variant
C1292780|T191|Therapy-Related Myelodysplastic Syndrome
C1292780|T191|Therapy Related Myelodysplastic Syndrome
C1292780|T191|Therapy-Related MDS
C1292780|T191|t-MDS
C1512738|T191|Infiltrating Bladder Urothelial Carcinoma, Lipid-Cell Variant
C0862432|T191|Stage IV Bladder Urothelial Carcinoma
C0862432|T191|Stage IV Transitional Cell Carcinoma of the Bladder
C0862432|T191|Stage IV Transitional Cell Carcinoma of the Urinary Bladder
C0862432|T191|Stage IV Bladder Urothelial Carcinoma AJCC v7
C0862432|T191|Stage IV Transitional Cell Carcinoma of Urinary Bladder
C0862432|T191|Stage IV Transitional Cell Carcinoma of Bladder
C0862432|T191|Stage IV Urinary Bladder Transitional Cell Carcinoma
C0747053|T061|Inguinal Orchiectomy
C0747053|T061|inguinal orchiectomy
C0279989|T191|Childhood Epithelioid Sarcoma
C0279989|T191|childhood epithelioid sarcoma
C0279989|T191|epithelioid sarcoma, childhood
C0279989|T191|pediatric epithelioid sarcoma
C0279989|T191|sarcoma, epithelioid, childhood
C0279989|T191|Pediatric Epithelioid Sarcoma
C0796563|T191|Localized Malignant Neoplasm
C0796563|T191|Localized Cancer
C0796563|T191|Localized Malignancy
C0796563|T191|local cancer
C0796563|T191|Local Cancer
C0278772|T191|Localized Resectable Adult Liver Carcinoma
C0278772|T191|liver cancer, localized resectable adult primary
C0278772|T191|Localized Resectable Adult Liver Cancer
C0278772|T191|hepatoma, localized resectable adult primary
C0278772|T191|adult primary liver cancer, localized resectable
C0278772|T191|Localized Resectable Adult Primary Cancer of the Liver
C0278772|T191|Localized Resectable Adult Primary Cancer of Liver
C0278772|T191|localized resectable adult primary liver cancer
C0278772|T191|Localized Resectable Adult Primary Liver Cancer
C0278772|T191|adult primary hepatoma, localized resectable
C3272446|T033|N1bI Stage Finding
C2698997|T191|Carcinoma Arising from Craniopharyngioma
C2698997|T191|CRANIOPHARYNGIOMA, MALIGNANT
C2698997|T191|CARCINOMA ARISING FROM CRANIOPHARYNGIOMA
C0027667|T191|Metastatic Malignant Neoplasm of Unknown Primary Origin
C0027667|T191|Metastatic Malignant Neoplasm of Unknown Primary
C0027667|T191|Metastatic Neoplasm of Unknown Primary Origin
C0027667|T191|Cancer of Unknown Primary Site
C0027667|T191|occult primary tumor
C0027667|T191|cancer of unknown primary origin
C2985170|T191|Multifocal Glioblastomas
C0280183|T191|Recurrent Grade 2 Follicular Lymphoma
C0280183|T191|Relapsed Grade II Follicular Mixed Cell Lymphoma
C0280183|T191|relapsed follicular mixed cell lymphoma
C0280183|T191|Relapsed Follicular Mixed Cell Lymphoma
C0280183|T191|recurrent grade 2 follicular lymphoma
C0280183|T191|Recurrent Grade II Follicular Lymphoma
C0280183|T191|Recurrent Follicular Mixed Cell Lymphoma
C0280183|T191|follicular mixed cell lymphoma, recurrent
C0280183|T191|Recurrent Grade II Follicular Mixed Cell Lymphoma
C0280183|T191|recurrent grade II follicular mixed cell lymphoma
C0280183|T191|follicular mixed cell lymphoma, relapsed
C0280183|T191|Relapsed Grade II Follicular Lymphoma
C0854776|T191|Unresectable Pancreatic Cancer
C0854776|T191|Non-Resectable Pancreatic Carcinoma
C0854776|T191|Pancreatic Carcinoma, Non-Resectable
C0854776|T191|Non-Resectable Pancreas Carcinoma
C0854776|T191|Unresectable Pancreatic Carcinoma
C0854776|T191|Non-Resectable Carcinoma of Pancreas
C0854776|T191|Non-Resectable Carcinoma of the Pancreas
C0854776|T191|Pancreatic carcinoma non-resectable
C1332287|T191|Anaplastic Malignant Neoplasm
C2986684|T191|Stage II AIDS-Related Lymphoma
C2986684|T191|stage II AIDS-related lymphoma
CL378319|T061|Intracavitary Balloon Brachytherapy
CL378319|T061|intracavitary balloon brachytherapy
C1334755|T191|Microinvasive Malignant Neoplasm
C0347019|T191|Metastatic Malignant Neoplasm to the Eye
C0347019|T191|Metastatic Neoplasm to the Eye
C0347019|T191|Eye Metastasis
C0347019|T191|Metastasis to the Eye
C0347019|T191|Metastasis to Eye
C0347019|T191|Metastatic Tumor to the Eye
C0347019|T191|Metastases to Eye
C0347019|T191|Metastases to the Eye
C1512751|T191|Infiltrating Urothelial Carcinoma
C1512751|T191|Infiltrating Transitional Cell Carcinoma of the Urinary Tract
C0279646|T191|Childhood Acute Monocytic Leukemia
C0279646|T191|childhood acute monocytic leukemia with differentiation
C0279646|T191|pediatric acute monocytic leukemia
C0279646|T191|Pediatric Acute Differentiated Monocytic Leukemia
C0279646|T191|pediatric AMOL, differentiated
C0279646|T191|childhood AMOL
C0279646|T191|monocytic leukemia with differentiation, childhood acute
C0279646|T191|childhood AMOL, differentiated
C0279646|T191|AMOL, childhood
C0279646|T191|acute monocytic leukemia, childhood
C0279646|T191|childhood acute monocytic leukemia (M5b)
C0279646|T191|M5b childhood acute monocytic leukemia with differentiation
C0279646|T191|acute monocytic leukemia with differentiation, childhood
C0279646|T191|childhood acute M5b leukemia
C0279646|T191|M5b childhood AMOL, differentiated
C0279646|T191|Childhood Acute M5b Leukemia
C0279646|T191|M5b Pediatric Acute Differentiated Monocytic Leukemia
C0279646|T191|Childhood Acute Monocytic Leukemia with Differentiation
C0279646|T191|Pediatric Acute M5b Leukemia
C0279646|T191|childhood acute differentiated monocytic leukemia (M5b)
C0279646|T191|AMOL, pediatric
C0279646|T191|pediatric AMOL
C0279646|T191|pediatric acute monocytic leukemia with differentiation
C0279646|T191|leukemia, childhood acute monocytic
C0279646|T191|pediatric acute M5b leukemia
C0279646|T191|Pediatric Acute Monocytic Leukemia with Differentiation
C0279646|T191|M5b leukemia, childhood acute
C0279646|T191|M5b Childhood Acute Differentiated Monocytic Leukemia
C0279646|T191|leukemia, childhood acute monocytic with differentiation
C0279646|T191|pediatric acute differentiated monocytic leukemia
C0279646|T191|monocytic leukemia, childhood acute
C0279646|T191|Childhood Acute Differentiated Monocytic Leukemia (M5b)
C0279646|T191|M5b pediatric acute monocytic leukemia with differentiation
C0854198|T191|Metastatic Malignant Neoplasm to the Abdominal Cavity
C0854198|T191|Metastatic Neoplasm to the Abdominal Cavity
C0854198|T191|Metastatic Tumor to the Abdominal Cavity
C0854198|T191|Metastases to the Abdominal Cavity
C0854198|T191|Metastasis to the Abdominal Cavity
CL416259|T191|Secondary Central Nervous System Hodgkin Lymphoma
CL416259|T191|secondary central nervous system Hodgkin lymphoma
C1334272|T191|Invasive Apocrine Breast Carcinoma
C1334272|T191|Infiltrating Apocrine Carcinoma of the Breast
C1334272|T191|Invasive Apocrine Carcinoma of the Breast
C1334272|T191|Infiltrating Apocrine Breast Carcinoma
C1334272|T191|Invasive Apocrine Carcinoma of Breast
C1334272|T191|Infiltrating Apocrine Carcinoma of Breast
C1720728|T191|AIDS Related Immunoblastic Lymphoma
C1720728|T191|AIDS-related immunoblastic large cell lymphoma
C1720728|T191|immunoblastic large cell lymphoma, AIDS-related
C1720728|T191|AIDS Related Immunoblastic Large Cell Lymphoma
C1720728|T191|Immunoblastic sarcoma associated with AIDS
C1720728|T191|Immunoblastic lymphoma associated with AIDS
C1720728|T191|AIDS-Associated Immunoblastic Large Cell Lymphoma
C1720728|T191|AIDS-associated immunoblastic large cell lymphoma
C1720728|T191|Immunoblastic lymphoma associated with AIDS (disorder)
C1720728|T191|AIDS Associated Immunoblastic Lymphoma
C115204|T191|Childhood Grade III Lymphomatoid Granulomatosis
C0280240|T191|Localized Urothelial Carcinoma of the Renal Pelvis and Ureter
C0280240|T191|Localized Transitional Cell Cancer of Renal Pelvis and Ureter
C0280240|T191|Localized Transitional Cell Cancer of the Renal Pelvis and Ureter
C0280240|T191|Localized Transitional Cell Carcinoma of Renal Pelvis and Ureter
C1332968|T191|Childhood Extraskeletal Osteosarcoma
C1332968|T191|Pediatric Extraosseous Osteosarcoma
C1332968|T191|Pediatric Extraskeletal Osteosarcoma
C1332968|T191|Childhood Extraosseous Osteosarcoma
C0279582|T191|Childhood Burkitt Leukemia
C0279582|T191|leukemia, childhood acute lymphocytic , L3
C0279582|T191|L3 acute lymphoblastic leukemia, childhood
C0279582|T191|L3 Childhood ALL
C0279582|T191|L3 Pediatric Acute Lymphocytic Leukemia
C0279582|T191|L3 childhood acute lymphoblastic leukemia
C0279582|T191|Pediatric Burkitt's Leukemia
C0279582|T191|L3 lymphoblastic leukemia, acute childhood
C0279582|T191|L3 childhood acute lymphocytic leukemia
C0279582|T191|childhood acute lymphoblastic leukemia, L3
C0279582|T191|pediatric ALL, L3
C0279582|T191|L3 pediatric ALL
C0279582|T191|L3 Pediatric Acute Lymphoblastic Leukemia
C0279582|T191|acute lymphoblastic leukemia, childhood L3
C0279582|T191|pediatric Burkitt's leukemia
C0279582|T191|childhood ALL, L3
C0279582|T191|pediatric acute lymphocytic leukemia, L3
C0279582|T191|ALL, L3 pediatric
C0279582|T191|acute lymphocytic leukemia, childhood L3
C0279582|T191|L3 Childhood Acute Lymphoblastic Leukemia
C0279582|T191|L3 acute lymphocytic leukemia, childhood
C0279582|T191|childhood acute lymphocytic leukemia, L3
C0279582|T191|pediatric acute lymphoblastic leukemia, L3
C0279582|T191|L3 Childhood Acute Lymphocytic Leukemia
C0279582|T191|ALL, pediatric L3
C0279582|T191|ALL, childhood L3
C0279582|T191|Childhood Burkitt's Leukemia
C0279582|T191|L3 Pediatric ALL
C0279582|T191|L3 lymphocytic leukemia, acute childhood
C0279582|T191|ALL, L3 childhood
C0279756|T034|Estrogen Receptor Negative
C0279756|T034|ER-
C0279756|T034|estrogen receptor negative
C0279756|T034|Negative Estrogen Receptor
C0279756|T034|negative estrogen receptor
C1335492|T191|Primary Systemic Anaplastic Large Cell Lymphoma, ALK-Positive
C1335492|T191|Primary Systemic ALK-Positive Anaplastic Large Cell Lymphoma
C1335492|T191|Primary Systemic ALK-Positive ALCL
C1335492|T191|Primary Systemic ALKoma
C3272451|T033|N1bIV Stage Finding
C0346300|T191|Pituitary Gland Carcinoma
C0346300|T191|Pituitary carcinoma (morphologic abnormality)
C0346300|T191|Carcinoma of the Pituitary Gland
C0346300|T191|Carcinoma of Pituitary Gland
C0346300|T191|Pituitary Cancer
C0346300|T191|Cancer of the Pituitary
C0346300|T191|Cancer of Pituitary Gland
C0346300|T191|Cancers, Pituitary
C0346300|T191|Pituitary gland cancer, NOS
C0346300|T191|Pituitary Cancers
C0346300|T191|Pituitary Gland Cancer
C0346300|T191|Cancer, Pituitary
C0346300|T191|Pituitary Carcinomas
C0346300|T191|Pituitary carcinoma, NOS
C0346300|T191|Cancer of the Pituitary Gland
C0346300|T191|Cancer of Pituitary
C0346300|T191|Carcinoma, Pituitary
C0346300|T191|Pituitary carcinoma (disorder)
C0346300|T191|Carcinoma of Pituitary
C0346300|T191|pituitary cancer
C0346300|T191|Pituitary Carcinoma
C0346300|T191|pituitary carcinoma
C0346300|T191|Carcinomas, Pituitary
C0346300|T191|Carcinoma of the Pituitary
C0346300|T191|Pituitary Gland Adenocarcinoma
C0346300|T191|Pituitary carcinoma
C0279584|T191|Childhood B Acute Lymphoblastic Leukemia
C0279584|T191|B-Cell Pediatric Acute Lymphoblastic Leukemia
C0279584|T191|Childhood Precursor B-Lymphoblastic Leukemia
C0279584|T191|B-Cell Childhood Acute Lymphogenous Leukemia
C0279584|T191|B Cell Pediatric Acute Lymphocytic Leukemia
C0279584|T191|B-Cell Pediatric Acute Lymphoid Leukemia
C0279584|T191|B-Cell Pediatric Acute Lymphogenous Leukemia
C0279584|T191|B-Cell Childhood Acute Lymphoid Leukemia
C0279584|T191|B-Cell Pediatric ALL
C0279584|T191|B Cell Childhood Acute Lymphocytic Leukemia
C0279584|T191|B-Cell Childhood ALL
C0279584|T191|B Cell Pediatric ALL
C0279584|T191|B-Cell Childhood Acute Lymphocytic Leukemia
C0279584|T191|B Cell Pediatric Acute Lymphoblastic Leukemia
C0279584|T191|B-Cell Childhood Acute Lymphoblastic Leukemia
C0279584|T191|B Cell Childhood Acute Lymphoblastic Leukemia
C0279584|T191|B Cell Childhood ALL
C0279584|T191|B-Cell Pediatric Acute Lymphocytic Leukemia
C1519481|T049|Sporadic Breast Tumor Mutation
C1519481|T049|Mutation in Sporadic Breast Tumor
C0278754|T191|Childhood Central Nervous System Germ Cell Tumor
C0278754|T191|Pediatric CNS Germ Cell Tumor
C0278754|T191|childhood germ cell CNS tumor
C0278754|T191|Childhood Germ Cell Neoplasm of the Central Nervous System
C0278754|T191|Childhood Germ Cell Tumor of CNS
C0278754|T191|Pediatric Germ Cell Tumor of the Central Nervous System
C0278754|T191|childhood CNS tumor, germ cell
C0278754|T191|Childhood Germ Cell Neoplasm of the CNS
C0278754|T191|childhood central nervous system germ cell tumor
C0278754|T191|Pediatric Germ Cell Tumor of Central Nervous System
C0278754|T191|Childhood Central Nervous System Germ Cell Neoplasm
C0278754|T191|Childhood Germ Cell Tumor of the CNS
C0278754|T191|Pediatric Germ Cell Neoplasm of the Central Nervous System
C0278754|T191|Pediatric Germ Cell Tumor of the CNS
C0278754|T191|Pediatric Germ Cell Neoplasm of Central Nervous System
C0278754|T191|Childhood Germ Cell Tumor of Central Nervous System
C0278754|T191|Pediatric Central Nervous System Germ Cell Neoplasm
C0278754|T191|central nervous system tumor, germ cell, childhood
C0278754|T191|childhood CNS germ cell tumor
C0278754|T191|Pediatric Germ Cell Neoplasm of CNS
C0278754|T191|Pediatric CNS Germ Cell Neoplasm
C0278754|T191|CNS tumor, childhood germ cell
C0278754|T191|Childhood Germ Cell Tumor of the Central Nervous System
C0278754|T191|Pediatric Germ Cell Neoplasm of the CNS
C0278754|T191|Childhood CNS Germ Cell Tumor
C0278754|T191|CNS tumor, pediatric germ cell
C0278754|T191|Childhood CNS Germ Cell Neoplasm
C0278754|T191|Childhood Germ Cell Neoplasm of CNS
C0278754|T191|Pediatric Central Nervous System Germ Cell Tumor
C0278754|T191|Childhood Germ Cell Neoplasm of Central Nervous System
C0278754|T191|Pediatric Germ Cell Tumor of CNS
C0278754|T191|germ cell CNS tumor, childhood
C0334224|T191|Malignant Neoplasm, Uncertain Whether Primary or Metastatic
C1708717|T191|Localized Resectable Adult Hepatocellular Carcinoma
C0854788|T191|Recurrent Small Intestinal Carcinoma
C0854788|T191|Recurrent Small Bowel Carcinoma
C0854788|T191|Relapsed Carcinoma of the Small Bowel
C0854788|T191|Recurrent Carcinoma of the Small Bowel
C0854788|T191|Recurrent Cancer of the Small Intestine
C0854788|T191|Relapsed Small Intestine Carcinoma
C0854788|T191|Relapsed Carcinoma of Small Bowel
C0854788|T191|Relapsed Small Intestine Cancer
C0854788|T191|Small intestine carcinoma recurrent
C0854788|T191|Small Intestine Carcinoma, Recurrent
C0854788|T191|recurrent small intestine cancer
C0854788|T191|small intestine cancer, recurrent
C0854788|T191|Recurrent Carcinoma of Small Bowel
C0854788|T191|Relapsed Carcinoma of Small Intestine
C0854788|T191|Relapsed Small Bowel Carcinoma
C0854788|T191|Relapsed Cancer of the Small Intestine
C0854788|T191|recurrent small bowel cancer
C0854788|T191|Recurrent Small Intestinal Cancer
C0854788|T191|Recurrent Carcinoma of the Small Intestine
C0854788|T191|small bowel cancer, recurrent
C0854788|T191|Recurrent Cancer of Small Intestine
C0854788|T191|Relapsed Carcinoma of the Small Intestine
C0854788|T191|Relapsed Cancer of Small Intestine
C0854788|T191|Recurrent Carcinoma of Small Intestine
C0854788|T191|Recurrent Small Intestine Carcinoma
C0851344|T110|Exemestane
C0851344|T110|FCE-24304
C0851344|T110|6-Methyleneandrosta-1,4-diene-3,17-dione
C0851344|T110|EXEMESTANE
C0851344|T110|Aromasin
C0851344|T110|exemestane
C1334149|T191|Iatrogenic Kaposi Sarcoma
C1334149|T191|Iatrogenic Kaposi's Sarcoma
C1335924|T191|Thymic Sarcomatoid Carcinoma
C1335924|T191|Thymic Carcinosarcoma
C1335924|T191|Sarcomatoid Carcinoma of the Thymus
C1335924|T191|Thymus Sarcomatoid Carcinoma
C1335924|T191|Sarcomatoid Carcinoma of Thymus
C1335924|T191|Thymic Spindle Cell Carcinoma
C1332899|T191|Cerebellar Glioblastoma
C1332899|T191|Grade IV Cerebellar Astrocytic Tumor
C1332899|T191|Cerebellar Glioblastoma Multiforme
C1332899|T191|Grade IV Astrocytic Neoplasm of the Cerebellum
C1332899|T191|Grade IV Astrocytic Tumor of the Cerebellum
C1332899|T191|Grade IV Astrocytic Neoplasm of Cerebellum
C1332899|T191|Glioblastoma of Cerebellum
C1332899|T191|Glioblastoma of the Cerebellum
C1332899|T191|Grade IV Astrocytic Tumor of Cerebellum
C1332899|T191|Grade IV Cerebellar Astrocytic Neoplasm
C0751483|T191|Hereditary Retinoblastoma
C0751483|T191|Familial Retinoblastoma
C0751483|T191|Retinoblastoma, Hereditary
C0751483|T191|Familial Retinoblastomas
C0751483|T191|hereditary retinoblastoma
C0751483|T191|Retinoblastomas, Hereditary
C0751483|T191|Hereditary Retinoblastomas
C0751483|T191|Retinoblastoma, Familial
C0751483|T191|Retinoblastomas, Familial
C0751483|T191|retinoblastoma, hereditary
C0854743|T191|Stage 0 AIDS-Related Anal Canal Cancer
C0854743|T191|Stage 0 AIDS-Related Anal Canal Cancer AJCC v6
C0854743|T191|Stage 0 AIDS-Related Anal Canal Cancer AJCC v7
C0362051|T191|Malignant Neoplasm of Multiple Primary Sites
C1439275|T191|Disseminated Carcinoma
C1439275|T191|Disseminated carcinoma
C0481121|T037|Oral Contraceptive
C0481121|T037|OC
C0481121|T037|Oral contraceptive
C0481121|T037|The pill
C0481121|T037|Pill - oral contraception
C0481121|T037|Oral contraceptive drug
C0481121|T037|Oral contraceptives
C0481121|T037|oral contraceptive
C0481121|T037|Oral Contraceptives
C0481121|T037|Oral contraceptive preparation
C0481121|T037|Birth control pill
C0481121|T037|Oral contraceptive agent
C0481121|T037|birth control pills
C0481121|T037|Inhibition of ovulation
C0481121|T037|OC - Oral contraceptive
C0481121|T037|Oral contraceptive agent (substance)
C0481121|T037|Pill
C0481121|T037|CONTRACEPTIVE PILLS FOR BIRTH CONTROL
C0481121|T037|Contraceptive pills for bc
C0481121|T037|Oral contraceptive preparation (product)
C0481121|T037|Oral contraception
C0481121|T037|birth control pill
C0481121|T037|Oral contraception (finding)
C0481121|T037|Oral Contraceptives causing adverse effects in therapeutic use
C0481121|T037|Contraceptives, Oral
C0481121|T037|Oral contraceptives causing adverse effects in therapeutic use
C1334442|T191|Lung Carcinoma Metastatic to the Liver
C1333600|T191|Hereditary Malignant Neoplasm
C1333600|T191|Hereditary Cancer
C1333600|T191|Familial Malignant Neoplasm
C1333600|T191|familial cancer
C1333600|T191|Familial Cancer
C0347023|T191|Metastatic Malignant Neoplasm to the Thyroid Gland
C0347023|T191|Metastatic Malignant Tumor to the Thyroid
C0347023|T191|Secondary Malignant Tumor to the Thyroid Gland
C0347023|T191|Metastatic Malignant Tumor to the Thyroid Gland
C0347023|T191|Metastatic Tumor to the Thyroid Gland
C0347023|T191|Secondary Malignant Tumor to the Thyroid
C0347023|T191|Metastasis to the Thyroid Gland
C0347023|T191|Metastatic Tumor to the Thyroid
C0347023|T191|Metastatic Malignant Neoplasm to the Thyroid
C0347023|T191|Secondary Malignant Neoplasm to the Thyroid
C0347023|T191|Metastatic Neoplasm to the Thyroid Gland
C0347023|T191|Metastasis to the Thyroid
C0347023|T191|Metastatic Neoplasm to the Thyroid
C0347023|T191|Secondary Malignant Neoplasm to the Thyroid Gland
C1335506|T191|Prostate Carcinoma Metastatic to the Lung
C0521174|T046|Microcalcification
C0521174|T046|Microcalcifications of the breast
C0521174|T046|microcalcifications
C0521174|T046|Microcalcification, calcified structure
C0521174|T046|Microcalcification, calcified structure (morphologic abnormality)
C0521174|T046|Microcalcifications of the breast (disorder)
C0521174|T046|microcalcification
C0521174|T046|Microcalcifications
C0521174|T046|Breast microcalcification
C0542407|T061|Total Abdominal Hysterectomy with Bilateral Salpingo-Oophorectomy
C1336815|T191|Transplant-Related Renal Cell Carcinoma
C0746341|T191|Recurrent Hodgkin Lymphoma
C0746341|T191|Recurrent Hodgkin's Disease
C0746341|T191|Hodgkin's disease recurrent
C0746341|T191|Hodgkin's disease NOS recurrent
C0746341|T191|Recurrent Hodgkin's Lymphoma
C1335720|T191|Recurrent Primitive Neuroectodermal Tumor
C2825306|T191|Therapy-Related Leukemia
C2825306|T191|Therapy Related Leukemia
C1336079|T191|Squamous Cell Breast Carcinoma
C1336079|T191|Primary Squamous Cell Breast Carcinoma
C1336079|T191|Primary Squamous Cell Carcinoma of the Breast
C1336079|T191|SCC of Breast
C1336079|T191|SCC of the Breast
C1336079|T191|Squamous Carcinoma of Breast
C1336079|T191|Squamous Cell Carcinoma of the Breast
C1336079|T191|Squamous Breast Carcinoma
C1336079|T191|Squamous Carcinoma of the Breast
C1336079|T191|Squamous Cell Carcinoma of Breast
C1336079|T191|Primary Squamous Cell Carcinoma of Breast
C0332377|T033|Tumor stage TX
C0332377|T033|TX Tumor Stage
C0332377|T033|TX Cancer Stage Finding
C0332377|T033|TX Primary Tumor Finding
C0332377|T033|TX Stage
C0332377|T033|TX Stage Finding
C0332377|T033|Tumour stage TX
C0332377|T033|TX stage
C0332377|T033|TX category
C0332377|T033|TX Tumor Finding
C0332377|T033|TX Primary Tumor Stage Finding
C0332377|T033|TX
C0332377|T033|TX category (finding)
C0332377|T033|TX TNM Finding
C0332377|T033|Tumor Stage TX
C0405348|T060|Excisional Biopsy of Breast
C1378463|T191|Recurrent Hypopharyngeal Carcinoma
C1378463|T191|Relapsed Carcinoma of the Hypopharynx
C1378463|T191|hypopharynx cancer, recurrent
C1378463|T191|recurrent hypopharyngeal cancer
C1378463|T191|Relapsed Cancer of the Hypopharynx
C1378463|T191|Relapsed Cancer of Hypopharynx
C1378463|T191|Recurrent Cancer of the Hypopharynx
C1378463|T191|Relapsed Carcinoma of Hypopharynx
C1378463|T191|Recurrent Carcinoma of the Hypopharynx
C1378463|T191|Relapsed Hypopharynx Carcinoma
C1378463|T191|Recurrent Hypopharynx Carcinoma
C1378463|T191|Relapsed Hypopharyngeal Cancer
C1378463|T191|Recurrent Hypopharyngeal Cancer
C1378463|T191|hypopharyngeal cancer, recurrent
C1378463|T191|Recurrent Carcinoma of Hypopharynx
C1378463|T191|Relapsed Hypopharyngeal Carcinoma
C1378463|T191|Recurrent Cancer of Hypopharynx
C1708781|T191|Lung Sarcomatoid Carcinoma
C1332945|T191|Childhood Botryoid-Type Embryonal Rhabdomyosarcoma of the Vagina
C1332945|T191|Vaginal Childhood Sarcoma Botryoides
C1332945|T191|Childhood Sarcoma Botryoides of the Vagina
C1332945|T191|Vaginal Childhood Botryoid-Type Embryonal Rhabdomyosarcoma
C1705285|T049|Mutation Abnormality
C1705285|T049|Genetic Change
C1705285|T049|Genetic Alteration
C1705285|T049|mutation
C1705285|T049|Mutated
C1705285|T049|Mutation
C0278510|T191|Childhood Medulloblastoma
C0278510|T191|infratentorial PNET, pediatric
C0278510|T191|PNET, childhood cerebellar
C0278510|T191|Medulloblastoma, Childhood
C0278510|T191|PNET, infratentorial, childhood
C0278510|T191|PNET, cerebellar, childhood
C0278510|T191|primitive neuroectodermal tumor, childhood infratentorial
C0278510|T191|medulloblastoma, childhood
C0278510|T191|pediatric medulloblastoma
C0278510|T191|childhood infratentorial PNET
C0278510|T191|primitive neuroectodermal tumor, pediatric infratentorial
C0278510|T191|Medulloblastomas, Childhood
C0278510|T191|infratentorial primitive neuroectodermal tumor, pediatric
C0278510|T191|Childhood Medulloblastomas
C0278510|T191|cerebellar PNET, childhood
C0278510|T191|PNET, infratentorial, pediatric
C0278510|T191|pediatric cerebellar PNET
C0278510|T191|cerebellar primitive neuroectodermal tumor, childhood
C0278510|T191|primitive neuroectodermal tumor, childhood cerebellar
C0278510|T191|PNET, pediatric cerebellar
C0278510|T191|infratentorial, childhood, PNET
C0278510|T191|pediatric infratentorial primitive neuroectodermal tumor
C0278510|T191|medulloblastoma, pediatric
C0278510|T191|PNET, childhood infratentorial
C0278510|T191|primitive neuroectodermal tumor, pediatric cerebellar
C0278510|T191|pediatric cerebellar primitive neuroectodermal tumor
C0278510|T191|PNET, pediatric infratentorial
C0278510|T191|PNET, cerebellar, pediatric
C0278510|T191|infratentorial, pediatric, PNET
C0278510|T191|childhood cerebellar primitive neuroectodermal tumor
C0278510|T191|infratentorial primitive neuroectodermal tumor, childhood
C0278510|T191|pediatric infratentorial PNET
C0278510|T191|cerebellar, childhood, PNET
C0278510|T191|Pediatric Medulloblastoma
C0278510|T191|infratentorial PNET, childhood
C0278510|T191|childhood cerebellar PNET
C0278510|T191|Brain tumor, child: Medulloblastoma
C0278510|T191|cerebellar PNET, pediatric
C0278510|T191|cerebellar primitive neuroectodermal tumor, pediatric
C0278510|T191|childhood infratentorial primitive neuroectodermal tumor
C0278510|T191|childhood medulloblastoma
C0278510|T191|cerebellar, pediatric, PNET
C104989|T061|Retreatment of Progressive Local Disease with External Beam Radiation
C1300990|T201|Tumor size, largest metastasis, additional dimension
C1300990|T201|Tumor size, largest metastasis, additional dimension (observable entity)
C1300990|T201|Tumour size, largest metastasis, additional dimension
C0030186|T191|Extramammary Paget Disease
C0030186|T191|PAGET DISEASE, EXTRAMAMMARY
C0030186|T191|Paget's disease, extramammary (except Paget's disease of bone) (morphologic abnormality)
C0030186|T191|Paget Disease, Extramammary [Disease/Finding]
C0030186|T191|Extramammary, Paget Disease
C0030186|T191|PAGET DIS EXTRA MAMMARY
C0030186|T191|Paget Disease, Extra-Mammary
C0030186|T191|Extramammary Paget's Disease
C0030186|T191|Paget's disease, extramammary (except Paget's disease of bone)
C0030186|T191|EXTRA MAMMARY PAGET DIS
C0030186|T191|Paget's Disease of the Skin
C0030186|T191|[M]Paget's disease, extramammary, excluding Paget's disease of bone
C0030186|T191|Paget disease, extramammary
C0030186|T191|Paget's Disease, Extra Mammary
C0030186|T191|PAGETS DIS EXTRAMAMMARY
C0030186|T191|Pagets Disease, Extramammary
C0030186|T191|Paget's Disease, Extra-Mammary
C0030186|T191|Extra-Mammary Paget Disease
C0030186|T191|Extra-Mammary Paget's Disease
C0030186|T191|Cutaneous Paget's Disease
C0030186|T191|Pagets Disease, Extra-Mammary
C0030186|T191|Paget Disease, Extra Mammary
C0030186|T191|Paget Disease Extramammary
C0030186|T191|Extra-Mammary Pagets Disease
C0030186|T191|Paget Disease, Extramammary
C0030186|T191|Extramammary Pagets Disease
C0030186|T191|EXTRA MAMMARY PAGETS DIS
C0030186|T191|Paget disease of skin
C0030186|T191|Paget's disease of skin
C0030186|T191|Extramammary Paget's disease
C0030186|T191|EXTRAMAMMARY PAGET DIS
C0030186|T191|Paget's Disease of Skin
C0030186|T191|PAGETS DIS EXTRA MAMMARY
C0030186|T191|PAGET DIS EXTRAMAMMARY
C0030186|T191|EXTRAMAMMARY PAGETS DIS
C0030186|T191|Extra Mammary Paget Disease
C0030186|T191|Paget's disease of skin (morphologic abnormality)
C0030186|T191|Paget's Disease, Extramammary
C0030186|T191|Extra Mammary Paget's Disease
C0030186|T191|Paget disease, extramammary (except Paget disease of bone)
C0030186|T191|Paget's Skin Disease
C1709094|T049|Transversion Mutation
C1709094|T049|Transversion
C1709094|T049|Nucleotide Transversion Abnormality
C1709094|T049|Multiple Transversion Mutations
C1709094|T049|transversion mutation
C1709094|T049|Mutation, Transversion
C1709094|T049|Transversion Mutations
C1709094|T049|Multiple Transversion Abnormalities
C1709448|T033|Painful Mass
C0445079|T033|N2a Stage Finding
C0445079|T033|N2a Lymph Node Finding
C0445079|T033|Lymph Node Stage N2a
C0445079|T033|Node stage N2a (finding)
C0445079|T033|N2a Stage
C0445079|T033|N2a Regional Lymph Nodes Finding
C0445079|T033|Node Stage N2a
C0445079|T033|N2a
C0445079|T033|N2a Node Finding
C0445079|T033|Node stage N2a
C0445079|T033|N2a Lymph Node Stage
C0445079|T033|N2a Cancer Stage Finding
C0445079|T033|N2a Node Stage
C0445079|T033|N2a TNM Finding
C0445079|T033|N2a Regional Lymph Node Stage Finding
C0854745|T191|Stage II AIDS-Related Anal Canal Cancer
C0854745|T191|Stage II AIDS-Related Anal Canal Cancer AJCC v6
C0854745|T191|Stage II AIDS-Related Anal Canal Cancer AJCC v7
C0279612|T191|Childhood Embryonal Rhabdomyosarcoma
C0279612|T191|embryonal childhood rhabdomyosarcoma
C0279612|T191|rhabdomyosarcoma, embryonal childhood
C0279612|T191|rhabdomyosarcoma, childhood embryonal
C0279612|T191|embryonal pediatric rhabdomyosarcoma
C0279612|T191|Pediatric Embryonal Rhabdomyosarcoma
C0279612|T191|pediatric rhabdomyosarcoma, embryonal
C0279612|T191|Embryonal Childhood Rhabdomyosarcoma
C0279612|T191|rhabdomyosarcoma, pediatric embryonal
C0279612|T191|childhood rhabdomyosarcoma, embryonal
C3272457|T033|N1mi Stage Finding
C1332274|T191|Paget Disease of the Anus
C1332274|T191|Paget's Disease of Anus
C1332274|T191|Anal Paget's Disease
C1332274|T191|Paget's Disease of the Anus
C1302660|T201|Secondary tumor size
C1302660|T201|Secondary tumour size
C1302660|T201|Secondary tumor size (observable entity)
C0024883|T061|Modified Radical Mastectomy
C0024883|T061|Mastectomies, Modified
C0024883|T061|Radical Mastectomies, Modified
C0024883|T061|MODIFIED RADICAL MASTECTOMY
C0024883|T061|Radical Mastectomy, Modified
C0024883|T061|Modified Mastectomy
C0024883|T061|Mastectomies, Modified Radical
C0024883|T061|Mastectomy, Modified
C0024883|T061|Modified Mastectomies
C0024883|T061|modified radical mastectomy
C0024883|T061|Modified radical mastectomy
C0024883|T061|Modified Radical Mastectomies
C0024883|T061|Modified radical mastectomy (procedure)
C0024883|T061|Mastectomy, Modified Radical
C1511542|T201|Craniospinal Axis Irradiation in Children
C1879494|T061|A-T-C Regimen
C1879494|T061|Adriamycin-Taxol-Cytoxan Regimen
C0278502|T191|Recurrent Gastric Carcinoma
C0278502|T191|Recurrent Cancer of Stomach
C0278502|T191|Stomach carcinoma recurrent
C0278502|T191|Recurrent Carcinoma of the Stomach
C0278502|T191|Recurrent Stomach Carcinoma
C0278502|T191|Recurrent Carcinoma of Stomach
C0278502|T191|Recurrent Gastric Cancer
C0278502|T191|stomach cancer, recurrent
C0278502|T191|Stomach cancer recurrent
C0278502|T191|Gastric cancer recurrent
C0278502|T191|Gastric carcinoma recurrent
C0278502|T191|Gastric Carcinoma, Recurrent
C0278502|T191|gastric cancer, recurrent
C0278502|T191|Recurrent Stomach Cancer
C0278502|T191|Recurrent Cancer of the Stomach
C0278502|T191|recurrent gastric cancer
C0220647|T191|Carcinoma of Unknown Primary Origin
C0220647|T191|CUP
C0220647|T191|carcinoma of unknown primary
C0220647|T191|Carcinoma of Unknown Primary
C0281293|T191|AIDS-Related Hodgkin Lymphoma
C0281293|T191|HIV-Associated Hodgkin's Disease
C0281293|T191|HIV-Related Hodgkin's Disease
C0281293|T191|HIV-Related Hodgkin's Lymphoma
C0281293|T191|AIDS-Associated Hodgkin's Disease
C0281293|T191|AIDS-Related Hodgkin's Disease
C0281293|T191|AIDS-Related Hodgkin's Lymphoma
C0281293|T191|AIDS-Associated Hodgkin's Lymphoma
C0281293|T191|HIV-Associated Hodgkin's Lymphoma
C0281293|T191|AIDS-related Hodgkin lymphoma
C1514507|T191|Prostate Basal Cell Carcinoma
C1514507|T191|Basal Cell Carcinoma of the Prostate
C0475751|T033|Tumor stage T4
C0475751|T033|T4 Tumor Finding
C0475751|T033|Tumour stage T4
C0475751|T033|T4 category
C0475751|T033|T4 category (finding)
C0475751|T033|T4 Stage Finding
C0475751|T033|T4 Stage
C0475751|T033|T4 tumor stage
C0475751|T033|T4 Primary Tumor Stage Finding
C0475751|T033|T4 TNM Finding
C0475751|T033|T4
C0475751|T033|T4 Cancer Stage Finding
C0475751|T033|T4 Tumor Stage
C0475751|T033|T4 stage
C0475751|T033|T4 Primary Tumor Finding
C0475751|T033|Tumor Stage T4
C1831735|T061|Tomotherapy
C1831735|T061|Helical Tomotherapy
C1831735|T061|tomotherapy
C1831735|T061|Tomotherapy, Helical
C1831735|T061|helical tomotherapy
C1831735|T061|Helical Tomotherapies
C1831735|T061|Tomotherapies, Helical
C1334792|T191|Moderately Differentiated Prostate Adenocarcinoma
C0596611|T045|Gene Mutation
C0596611|T045|Gene mutation
C0596611|T045|Sequence Alteration
C0596611|T045|Gene Alteration
C0596611|T045|MOLPATH.MUT
C0596611|T045|DNA Sequence Alteration
C0596611|T045|DNA Alteration
C0596611|T045|gene mutation
C0475412|T082|Goiter size
C0475412|T082|Goitre size
C0475412|T082|Size of goitre
C0475412|T082|Size of goiter
C0475412|T082|Goiter size (observable entity)
C0280483|T191|Adult Anaplastic Astrocytoma
C0280483|T191|Adult Grade III Astrocytoma
C0280483|T191|Undifferentiated Astrocytoma of Adult
C0280483|T191|astrocytoma, adult anaplastic
C0280483|T191|Undifferentiated Astrocytoma of the Adult
C0280483|T191|Grade III Adult Astrocytic Neoplasm
C0280483|T191|Anaplastic Astrocytoma of the Adult
C0280483|T191|Grade III Adult Astrocytic Tumor
C0280483|T191|adult anaplastic astrocytoma
C0280483|T191|Grade III Adult Astrocytoma
C0280483|T191|Anaplastic Astrocytoma of Adult
C0280483|T191|anaplastic astrocytoma, adult
C0280483|T191|Adult Undifferentiated Astrocytoma
C1335694|T191|Recurrent Bone Ewing Sarcoma
C1335694|T191|Recurrent Osseous Ewing's Sarcoma
C1335694|T191|Relapsed Ewing's Sarcoma of Bone
C1335694|T191|Relapsed Osseous Ewing's Sarcoma
C1335694|T191|Recurrent Ewing's Sarcoma of Bone
C1335694|T191|Relapsed Skeletal Ewing's Sarcoma
C1335694|T191|Relapsed Bone Ewing's Sarcoma
C1335694|T191|Relapsed Ewing's Sarcoma of the Bone
C1335694|T191|Recurrent Bone Ewing's Sarcoma
C1335694|T191|Recurrent Skeletal Ewing's Sarcoma
C1335694|T191|Recurrent Ewing's Sarcoma of the Bone
C0553989|T060|Excisional Biopsy of Lymph Node
C0553989|T060|Lymph Node Excision
C104919|T061|Cobalt-60 Radiation Therapy
C0278844|T191|Childhood Immunoblastic Lymphoma
C0278844|T191|Pediatric Immunoblastic Lymphoma
C0278844|T191|childhood immunoblastic large cell lymphoma
C0278844|T191|lymphoma, immunoblastic large cell childhood
C0278844|T191|immunoblastic large cell lymphoma, childhood
C0278844|T191|Childhood Immunoblastic Large Cell Lymphoma
C0278844|T191|pediatric IBL lymphoma
C0278844|T191|large cell lymphoma, childhood immunoblastic
C0278844|T191|IBL lymphoma, childhood
C0278844|T191|pediatric immunoblastic large cell lymphoma
C0278844|T191|Pediatric Immunoblastic Large Cell Lymphoma
C0278844|T191|childhood IBL lymphoma
C0279525|T191|Childhood Lymphoblastic Lymphoma
C0279525|T191|non-Hodgkin's lymphoma, childhood lymphoblastic
C0279525|T191|CLNHL
C0279525|T191|NHL, childhood lymphoblastic
C0279525|T191|lymphoma, childhood lymphoblastic non-Hodgkin's
C0279525|T191|pediatric lymphoblastic lymphoma
C0279525|T191|Childhood Precursor Lymphoblastic Lymphoma
C0279525|T191|lymphoblastic non-Hodgkin's lymphoma, childhood
C0279525|T191|lymphoblastic lymphoma, childhood
C0279525|T191|Pediatric Lymphoblastic Lymphoma
C0279525|T191|pediatric lymphoblastic non-Hodgkin's lymphoma
C0279525|T191|lymphoblastic lymphoma, pediatric
C0279525|T191|lymphoma, pediatric lymphoblastic
C0279525|T191|lymphoma, childhood lymphoblastic
C0279525|T191|childhood lymphoblastic lymphoma
C0860580|T191|Medullary Breast Carcinoma
C0860580|T191|ductal medullary breast carcinoma with lymphocytic infiltrate
C0860580|T191|Invasive Medullary Carcinoma of the Breast
C0860580|T191|Invasive Medullary Carcinoma of Breast
C0860580|T191|Medullary Breast Carcinoma with Lymphoid Stroma
C0860580|T191|Infiltrating Medullary Carcinoma of the Breast
C0860580|T191|Medullary Carcinoma of the Breast
C0860580|T191|Invasive Medullary Breast Carcinoma
C0860580|T191|medullary ductal breast carcinoma with lymphocytic infiltrate
C0860580|T191|Medullary Carcinoma of Breast
C0860580|T191|Infiltrating Medullary Carcinoma of Breast
C0860580|T191|medullary breast carcinoma
C0860580|T191|Medullary carcinoma of breast
C1377599|T191|Childhood Central Nervous System Teratoma
C1377599|T191|Pediatric Teratoma of Central Nervous System
C1377599|T191|Childhood Teratoma of CNS
C1377599|T191|Childhood CNS Teratoma
C1377599|T191|Pediatric Central Nervous System Teratoma
C1377599|T191|Childhood Teratoma of the CNS
C1377599|T191|Pediatric Teratoma of the Central Nervous System
C1377599|T191|Pediatric Teratoma of CNS
C1377599|T191|childhood central nervous system teratoma
C1377599|T191|Childhood Teratoma of Central Nervous System
C1377599|T191|Pediatric Teratoma of the CNS
C1377599|T191|Childhood Teratoma of the Central Nervous System
C1377599|T191|Pediatric CNS Teratoma
C1377599|T191|childhood CNS teratoma
C1332984|T191|Childhood Myxoid Chondrosarcoma
C1332984|T191|Pediatric Myxoid Chondrosarcoma
C1134719|T191|Invasive Ductal Carcinoma, Not Otherwise Specified
C1134719|T191|Invasive Ductal Carcinoma, No Specific Type
C1134719|T191|Invasive Ductal Breast Carcinoma
C1134719|T191|Infiltrating Ductal Carcinoma of the Breast
C1134719|T191|Infiltrating Ductal Carcinoma of Breast
C1134719|T191|Invasive Ductal Carcinoma of the Breast
C1134719|T191|Invasive Ductal Adenocarcinoma
C1134719|T191|Infiltrating Ductal Adenocarcinoma
C1134719|T191|Infiltrating Ductal Carcinoma
C1134719|T191|Invasive Ductal Carcinoma, NST
C1134719|T191|Invasive Ductal Carcinoma
C1134719|T191|Infiltrating Ductal Breast Carcinoma
C1134719|T191|Invasive Ductal Carcinoma, NOS
C1134719|T191|Invasive Ductal Carcinoma of Breast
C1134719|T191|infiltrating ductal carcinoma
C0855089|T191|Recurrent B-Cell Non-Hodgkin Lymphoma
C0855089|T191|B-Cell Lymphoma Recurrent
C0855089|T191|Recurrent B-Cell Lymphoma
C0855089|T191|Recurrent B-Cell Non-Hodgkin's Lymphoma
C0347001|T191|Metastatic Malignant Neoplasm to the Prostate
C0347001|T191|Metastasis to Prostate
C0347001|T191|Metastatic Tumor to the Prostate
C0347001|T191|Metastatic Neoplasm to the Prostate
C0347001|T191|Metastases to the Prostate
C0347001|T191|Metastasis to the Prostate
C0347001|T191|Metastases to Prostate
C1514587|T033|Pseudoencapsulated Mass
C1334791|T191|Moderately Differentiated Malignant Neoplasm
C0278517|T191|Recurrent Non-Small Cell Lung Carcinoma
C0278517|T191|Non Small Cell Lung Cancer, Recurrent
C0278517|T191|Recurrent Non-Small Cell Lung Cancer
C0278517|T191|Recurrent Non-Small Cell Cancer of the Lung
C0278517|T191|Recurrent Non-Small Cell Cancer of Lung
C0278517|T191|Recurrent NSCLC
C0278517|T191|Non Small Cell Lung Cancer Recurrent
C0854843|T191|Recurrent Enteropathy-Associated T-Cell Lymphoma
C0854843|T191|Relapsed Intestinal T-Cell Lymphoma
C0854843|T191|Recurrent Intestinal T-Cell Lymphoma
C0854843|T191|Recurrent Enteropathy-type T-Cell Lymphoma
C1332613|T191|Breast Adenocarcinoma with Squamous Metaplasia
C1332613|T191|Adenocarcinoma of the Breast with Squamous Metaplasia
C1332613|T191|Adenocarcinoma of Breast with Squamous Metaplasia
C1332613|T191|Adenoacanthoma of the Breast
C1332613|T191|Breast Adenoacanthoma
C1332613|T191|Adenoacanthoma of Breast
C0041687|T061|Unilateral Oophorectomy
C0041687|T061|Unilateral oophorectomy
C0041687|T061|ovariectomy - unilateral
C0041687|T061|Unilateral excision of ovary
C0041687|T061|Unilateral excision of ovary (situation)
C0041687|T061|Unilateral Ovariectomy
C0041687|T061|Oophorectomy unilateral
C0278727|T191|Recurrent Small Cell Lung Carcinoma
C0278727|T191|Recurrent Small Cell Carcinoma of Lung
C0278727|T191|small cell lung cancer, recurrent
C0278727|T191|oat cell lung cancer, recurrent
C0278727|T191|Relapsed Small Cell Lung Carcinoma
C0278727|T191|Relapsed Small Cell Lung Cancer
C0278727|T191|Small cell lung cancer recurrent
C0278727|T191|recurrent SCLC
C0278727|T191|lung cancer, recurrent small cell
C0278727|T191|SCLC, recurrent
C0278727|T191|Recurrent Small Cell Lung Cancer
C0278727|T191|Relapsed Small Cell Carcinoma of Lung
C0278727|T191|Recurrent Small Cell Carcinoma of the Lung
C0278727|T191|recurrent small cell lung cancer
C0278727|T191|Relapsed Small Cell Carcinoma of the Lung
C0280392|T191|Recurrent Hypopharyngeal Squamous Cell Carcinoma
C0280392|T191|recurrent squamous cell carcinoma of the hypopharynx
C0280392|T191|Recurrent Epidermoid Carcinoma of the Hypopharynx
C0280392|T191|hypopharyngeal squamous cell carcinoma, recurrent
C0280392|T191|Hypopharyngeal squamous cell carcinoma recurrent
C0280392|T191|Relapsed Squamous Cell Carcinoma of the Hypopharynx
C0280392|T191|Relapsed Hypopharyngeal Epidermoid Carcinoma
C0280392|T191|Recurrent Epidermoid Carcinoma of Hypopharynx
C0280392|T191|Relapsed Epidermoid Carcinoma of Hypopharynx
C0280392|T191|Recurrent Squamous Cell Carcinoma of Hypopharynx
C0280392|T191|hypopharynx squamous cell carcinoma, recurrent
C0280392|T191|Relapsed Epidermoid Carcinoma of the Hypopharynx
C0280392|T191|Recurrent Squamous Cell Carcinoma of the Hypopharynx
C0280392|T191|squamous cell carcinoma of the hypopharynx, recurrent
C0280392|T191|Relapsed Hypopharyngeal Squamous Cell Carcinoma
C0280392|T191|Recurrent Hypopharyngeal Epidermoid Carcinoma
C0280392|T191|epidermoid carcinoma of the hypopharynx, recurrent
C0280392|T191|Relapsed Squamous Cell Carcinoma of Hypopharynx
C0280392|T191|Squamous cell carcinoma of the hypopharynx recurrent
C0248241|T061|FEC Regimen
C0248241|T061|fluorouracil-epirubicin-cyclophosphamide Regimen
C0248241|T061|cyclophosphamide/epirubicin/fluorouracil
C0248241|T061|FEC 100
C0248241|T061|CEF regimen
C0248241|T061|CTX/EPI/5-FU
C0248241|T061|Fluorouracil-Epirubicin-Cytoxan Regimen
C0248241|T061|FEC
C0248241|T061|CEF Regimen
C0248241|T061|CEF
C0248241|T061|FEC regimen
C0248241|T061|FEC protocol
C0248241|T061|Cyclophosphamide/Epirubicin/Fluorouracil
C0855013|T191|Recurrent Chondrosarcoma
C0855013|T191|Relapsed Chondrosarcoma
C0855013|T191|Chondrosarcoma, Recurrent
C0855013|T191|Chondrosarcoma recurrent
C1275593|T201|Lesion size, largest dimension
C1275593|T201|Lesion size, greatest dimension
C1275593|T201|Lesion size, largest dimension (observable entity)
C1300585|T191|Prostate Small Cell Carcinoma
C1300585|T191|Oat Cell Carcinoma of the Prostate
C1300585|T191|Prostate Small Cell NEC
C1300585|T191|Small cell carcinoma of prostate (disorder)
C1300585|T191|Prostate Small Cell Neuroendocrine Carcinoma
C1300585|T191|Prostate Oat Cell Carcinoma
C1300585|T191|Oat Cell Carcinoma of Prostate
C1300585|T191|Small Cell Carcinoma of the Prostate
C1300585|T191|Small Cell Carcinoma of Prostate
C1300585|T191|Small cell carcinoma of prostate
C0441960|T033|N2 Stage Finding
C0441960|T033|N2 TNM Finding
C0441960|T033|N2 Stage
C0441960|T033|Node stage N2
C0441960|T033|N2 Cancer Stage Finding
C0441960|T033|Lymph Node Stage N2
C0441960|T033|N2
C0441960|T033|N2 Lymph Node Finding
C0441960|T033|N2 stage
C0441960|T033|Node Stage N2
C0441960|T033|N2 Regional Lymph Nodes Finding
C0441960|T033|N2 lymph node stage
C0441960|T033|N2 Node Stage
C0441960|T033|N2 Regional Lymph Node Stage Finding
C0441960|T033|N2 Node Finding
C0441960|T033|N2 category
C0441960|T033|N2 Lymph Node Stage
C0441960|T033|N2 category (finding)
C1711181|T033|Intraluminal Necrosis
C1332947|T191|Childhood Brain Anaplastic Astrocytoma
C1332947|T191|Grade III Childhood Brain Astrocytoma
C1332947|T191|Grade III Childhood Astrocytic Neoplasm of Brain
C1332947|T191|Grade III Pediatric Astrocytic Tumor of the Brain
C1332947|T191|Grade III Childhood Brain Astrocytic Tumor
C1332947|T191|Grade III Childhood Astrocytic Tumor of the Brain
C1332947|T191|Anaplastic Childhood Astrocytoma of the Brain
C1332947|T191|Anaplastic Pediatric Astrocytoma of Brain
C1332947|T191|Anaplastic Pediatric Brain Astrocytoma
C1332947|T191|Grade III Childhood Astrocytic Neoplasm of the Brain
C1332947|T191|Grade III Childhood Astrocytoma of Brain
C1332947|T191|Grade III Childhood Astrocytoma of the Brain
C1332947|T191|Grade III Pediatric Astrocytic Tumor of Brain
C1332947|T191|Grade III Pediatric Astrocytic Neoplasm of Brain
C1332947|T191|Grade III Pediatric Astrocytoma of Brain
C1332947|T191|Grade III Pediatric Astrocytoma of the Brain
C1332947|T191|Anaplastic Childhood Brain Astrocytoma
C1332947|T191|Grade III Pediatric Brain Astrocytoma
C1332947|T191|Grade III Pediatric Brain Astrocytic Tumor
C1332947|T191|Anaplastic Pediatric Astrocytoma of the Brain
C1332947|T191|Anaplastic Childhood Astrocytoma of Brain
C1332947|T191|Grade III Pediatric Brain Astrocytic Neoplasm
C1332947|T191|Grade III Childhood Astrocytic Tumor of Brain
C1332947|T191|Grade III Childhood Brain Astrocytic Neoplasm
C1332947|T191|Grade III Pediatric Astrocytic Neoplasm of the Brain
C1708263|T049|Guanosine to Thymidine Transversion Abnormality
C1708263|T049|Guanosine to Thymidine Mutation
C1708263|T049|Guanosine to Thymidine Transversion
C3273067|T191|Calcifying Nested Epithelial Stromal Tumor of the Liver
C0220611|T191|Childhood Rhabdomyosarcoma
C0220611|T191|childhood rhabdomyosarcoma
C0220611|T191|pediatric rhabdomyosarcoma
C0220611|T191|rhabdomyosarcoma, childhood
C0220611|T191|sarcoma, childhood rhabdomyosarcoma
C0220611|T191|Rhabdomyosarcoma, child
C0220611|T191|Pediatric Rhabdomyosarcoma
C0279649|T191|Childhood Acute Basophilic Leukemia
C0279649|T191|basophilic leukemia, childhood acute
C0279649|T191|pediatric acute basophilic leukemia
C0279649|T191|childhood acute basophilic leukemia
C0279649|T191|acute basophilic leukemia, childhood
C0279649|T191|leukemia, childhood acute basophilic
C0279649|T191|Pediatric Acute Basophilic Leukemia
C113812|T061|Involved-Field Radiation Therapy
C113812|T061|IFRT
C113812|T061|Involved field radiotherapy
C535972|T191|Lynch Syndrome
C535972|T191|Syndrome, Lynch
C535972|T191|COLORECTAL CANCER, HEREDITARY NONPOLYPOSIS, TYPE 1
C535972|T191|HNPCC - hereditary nonpolyposis colon cancer
C535972|T191|Lynch 1 Syndrome
C535972|T191|COLON CANCER, FAMILIAL NONPOLYPOSIS, TYPE 1
C535972|T191|Hereditary Nonpolyposis Colorectal Neoplasms
C535972|T191|HNPCC1
C535972|T191|Familial Non-Polyposis Colon Cancer Type 1
C535972|T191|Hereditary Non-Polyposis Colon Cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C535972|T191|Familial Non-Polyposis Colon Cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C535972|T191|Colorectal Neoplasms, Hereditary Nonpolyposis [Disease/Finding]
C535972|T191|Colon cancer, familial nonpolyposis, type 1
C535972|T191|hereditary colorectal endometrial cancer syndrome
C535972|T191|Lynch Cancer Family Syndrome I
C535972|T191|COLORECTAL NEOPL HEREDITARY NONPOLYPOSIS
C535972|T191|FCC1
C535972|T191|Hereditary nonpolyposis colon cancer (disorder)
C535972|T191|Lynch Syndrome I
C535972|T191|familial non-polyposis colon cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C535972|T191|Hereditary Non-Polyposis Colon Cancer
C535972|T191|Hereditary Nonpolyposis Colon Cancer
C535972|T191|LYNCH SYNDROME I
C535972|T191|hereditary non-polyposis colon cancer
C535972|T191|hereditary non-polyposis colon cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C535972|T191|Hereditary Nonpolyposis Colorectal Neoplasm
C535972|T191|HEREDITARY NONPOLYPOSIS COLORECTAL NEOPL
C535972|T191|COCA1
C535972|T191|Hereditary nonpolyposis colon cancer
C535972|T191|hereditary defective mismatch repair syndrome
C535972|T191|colon cancer, hereditary non-polyposis - Lynch syndrome
C535972|T191|Hereditary Defective Mismatch Repair Syndrome
C535972|T191|Colon Cancer, Familial Nonpolyposis
C535972|T191|hereditary nonpolyposis-Lynch syndrome
C535972|T191|Colorectal Cancer Hereditary Nonpolyposis
C535972|T191|Colorectal Neoplasms, Hereditary Nonpolyposis
C535972|T191|Hereditary Nonpolyposis Colorectal Cancer
C535972|T191|HNPCC
C535972|T191|hereditary nonpolyposis colon cancer
C535972|T191|Lynch syndrome
C535972|T191|Hereditary Non-Polyposis Colon Cancer Type 1
C535972|T191|Colorectal cancer, hereditary nonpolyposis, type 1
C535972|T191|Hereditary Colorectal Endometrial Cancer Syndrome
C0280186|T191|Recurrent Adult Burkitt Lymphoma
C0280186|T191|adult diffuse small cleaved cell lymphoma, relapsed
C0280186|T191|Recurrent Adult Burkitt's Lymphoma
C0280186|T191|Recurrent Adult Small Non-Cleaved Cell/Burkitt's Lymphoma
C0280186|T191|recurrent adult diffuse small cleaved cell lymphoma
C0280186|T191|small noncleaved cell lymphoma, recurrent, adult
C0280186|T191|Relapsed Adult Small Non-Cleaved Cell/Burkitt's Lymphoma
C0280186|T191|recurrent adult Burkitt lymphoma
C0280186|T191|adult diffuse small cleaved cell lymphoma, recurrent
C0280186|T191|relapsed adult small noncleaved cell lymphoma
C0280186|T191|diffuse small cleaved cell lymphoma, adult, recurrent
C0280186|T191|adult small noncleaved cell lymphoma, relapsed
C0280186|T191|small noncleaved cell lymphoma, adult, recurrent
C0280186|T191|recurrent adult diffuse small noncleaved cell/Burkitt's lymphoma
C0280186|T191|relapsed adult diffuse small cleaved cell lymphoma
C0280186|T191|Recurrent Adult Diffuse Small Non-Cleaved Cell Lymphoma
C0280186|T191|adult small noncleaved cell lymphoma, recurrent
C0280186|T191|diffuse small cleaved cell lymphoma, recurrent, adult
C0862601|T191|Vaginal Metastatic Adenocarcinoma
C0862601|T191|Vaginal adenocarcinoma metastatic
C0684817|T191|Metastatic Malignant Neoplasm to the Neck
C0684817|T191|Metastatic Neoplasm to the Neck
C0684817|T191|Metastases to Neck
C0684817|T191|Metastatic Tumor to the Neck
C0684817|T191|Metastasis to the Neck
C1333843|T191|Grade 3 Invasive Breast Carcinoma
C1333843|T191|Grade 3 Infiltrating Breast Carcinoma
C1333843|T191|Unfavorable Infiltrating Breast Carcinoma
C1333843|T191|Poorly Differentiated Infiltrating Breast Carcinoma
C1333843|T191|Poorly Differentiated Invasive Breast Carcinoma
C1333843|T191|High Combined Histologic Grade Infiltrating Breast Carcinoma
C0278684|T191|Recurrent Parathyroid Gland Carcinoma
C0278684|T191|Recurrent Parathyroid Carcinoma
C0278684|T191|Recurrent Parathyroid Cancer
C0278684|T191|carcinoma of the parathyroid, recurrent
C0278684|T191|cancer of the parathyroid, recurrent
C0278684|T191|recurrent parathyroid carcinoma
C0278684|T191|recurrent parathyroid cancer
C0278684|T191|parathyroid carcinoma, recurrent
C0278684|T191|parathyroid cancer, recurrent
